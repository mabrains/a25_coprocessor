module a25_coprocessor (i_clk,
    i_core_stall,
    i_fault,
    o_cache_enable,
    o_cache_flush,
    VPWR,
    VGND,
    i_copro_crm,
    i_copro_crn,
    i_copro_num,
    i_copro_opcode1,
    i_copro_opcode2,
    i_copro_operation,
    i_copro_write_data,
    i_fault_address,
    i_fault_status,
    o_cacheable_area,
    o_copro_read_data);
 input i_clk;
 input i_core_stall;
 input i_fault;
 output o_cache_enable;
 output o_cache_flush;
 input VPWR;
 input VGND;
 input [3:0] i_copro_crm;
 input [3:0] i_copro_crn;
 input [3:0] i_copro_num;
 input [2:0] i_copro_opcode1;
 input [2:0] i_copro_opcode2;
 input [1:0] i_copro_operation;
 input [31:0] i_copro_write_data;
 input [31:0] i_fault_address;
 input [7:0] i_fault_status;
 output [31:0] o_cacheable_area;
 output [31:0] o_copro_read_data;

 sky130_fd_sc_hd__clkbuf_2 _0507_ (.A(net53),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_2 _0508_ (.A(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(net53),
    .Y(_0173_));
 sky130_fd_sc_hd__buf_1 _0510_ (.A(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_2 _0511_ (.A(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(\disruptive_area[30] ),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(net7),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(net5),
    .Y(_0178_));
 sky130_fd_sc_hd__or4_4 _0515_ (.A(net8),
    .B(_0177_),
    .C(_0178_),
    .D(net6),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_2 _0516_ (.A(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__buf_2 _0517_ (.A(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_2 _0518_ (.A(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__buf_1 _0519_ (.A(net5),
    .X(_0183_));
 sky130_fd_sc_hd__or2_2 _0520_ (.A(net8),
    .B(net7),
    .X(_0184_));
 sky130_fd_sc_hd__or3_4 _0521_ (.A(_0183_),
    .B(net6),
    .C(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_4 _0522_ (.A(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(net120),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(net6),
    .Y(_0188_));
 sky130_fd_sc_hd__buf_1 _0525_ (.A(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__or3_4 _0526_ (.A(_0178_),
    .B(_0189_),
    .C(_0184_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_2 _0527_ (.A(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(\updateable_area[30] ),
    .Y(_0192_));
 sky130_fd_sc_hd__or4_4 _0529_ (.A(_0183_),
    .B(net6),
    .C(net8),
    .D(_0177_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_2 _0530_ (.A(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__or4_4 _0531_ (.A(_0178_),
    .B(_0189_),
    .C(net8),
    .D(_0177_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _0532_ (.A(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__or2b_1 _0533_ (.A(_0196_),
    .B_N(\fault_address[30] ),
    .X(_0197_));
 sky130_fd_sc_hd__o221a_1 _0534_ (.A1(_0187_),
    .A2(_0191_),
    .B1(_0192_),
    .B2(_0194_),
    .C1(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__o211ai_1 _0535_ (.A1(_0176_),
    .A2(_0182_),
    .B1(_0186_),
    .C1(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__a22o_1 _0536_ (.A1(net152),
    .A2(_0172_),
    .B1(_0175_),
    .B2(_0199_),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_2 _0537_ (.A(_0172_),
    .X(_0200_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\disruptive_area[29] ),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(net118),
    .Y(_0202_));
 sky130_fd_sc_hd__buf_2 _0540_ (.A(_0190_),
    .X(_0203_));
 sky130_fd_sc_hd__buf_2 _0541_ (.A(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(\fault_address[29] ),
    .Y(_0205_));
 sky130_fd_sc_hd__clkbuf_2 _0543_ (.A(_0195_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_2 _0544_ (.A(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(\updateable_area[29] ),
    .Y(_0208_));
 sky130_fd_sc_hd__buf_2 _0546_ (.A(_0193_),
    .X(_0209_));
 sky130_fd_sc_hd__o22a_1 _0547_ (.A1(_0205_),
    .A2(_0207_),
    .B1(_0208_),
    .B2(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__o221ai_1 _0548_ (.A1(_0201_),
    .A2(_0182_),
    .B1(_0202_),
    .B2(_0204_),
    .C1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__a22o_1 _0549_ (.A1(_0200_),
    .A2(net150),
    .B1(_0175_),
    .B2(_0211_),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(\disruptive_area[28] ),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(net117),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _0552_ (.A(\fault_address[28] ),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(\updateable_area[28] ),
    .Y(_0215_));
 sky130_fd_sc_hd__clkbuf_2 _0554_ (.A(_0194_),
    .X(_0216_));
 sky130_fd_sc_hd__o22a_1 _0555_ (.A1(_0214_),
    .A2(_0207_),
    .B1(_0215_),
    .B2(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__o221ai_2 _0556_ (.A1(_0212_),
    .A2(_0182_),
    .B1(_0213_),
    .B2(_0204_),
    .C1(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__a22o_1 _0557_ (.A1(_0200_),
    .A2(net149),
    .B1(_0175_),
    .B2(_0218_),
    .X(_0167_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(\disruptive_area[27] ),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(net116),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _0560_ (.A(\fault_address[27] ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(\updateable_area[27] ),
    .Y(_0222_));
 sky130_fd_sc_hd__o22a_1 _0562_ (.A1(_0221_),
    .A2(_0207_),
    .B1(_0222_),
    .B2(_0216_),
    .X(_0223_));
 sky130_fd_sc_hd__o221ai_1 _0563_ (.A1(_0219_),
    .A2(_0182_),
    .B1(_0220_),
    .B2(_0204_),
    .C1(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__a22o_1 _0564_ (.A1(_0200_),
    .A2(net148),
    .B1(_0175_),
    .B2(_0224_),
    .X(_0166_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(\disruptive_area[26] ),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(net115),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(\fault_address[26] ),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(\updateable_area[26] ),
    .Y(_0228_));
 sky130_fd_sc_hd__o22a_1 _0569_ (.A1(_0227_),
    .A2(_0207_),
    .B1(_0228_),
    .B2(_0216_),
    .X(_0229_));
 sky130_fd_sc_hd__o221ai_2 _0570_ (.A1(_0225_),
    .A2(_0182_),
    .B1(_0226_),
    .B2(_0204_),
    .C1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__a22o_1 _0571_ (.A1(_0200_),
    .A2(net147),
    .B1(_0175_),
    .B2(_0230_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _0572_ (.A(_0174_),
    .X(_0231_));
 sky130_fd_sc_hd__inv_2 _0573_ (.A(\disruptive_area[25] ),
    .Y(_0232_));
 sky130_fd_sc_hd__buf_4 _0574_ (.A(_0180_),
    .X(_0233_));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(net114),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0576_ (.A(\fault_address[25] ),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(\updateable_area[25] ),
    .Y(_0236_));
 sky130_fd_sc_hd__o22a_1 _0578_ (.A1(_0235_),
    .A2(_0207_),
    .B1(_0236_),
    .B2(_0216_),
    .X(_0237_));
 sky130_fd_sc_hd__o221ai_2 _0579_ (.A1(_0232_),
    .A2(_0233_),
    .B1(_0234_),
    .B2(_0204_),
    .C1(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__a22o_1 _0580_ (.A1(_0200_),
    .A2(net146),
    .B1(_0231_),
    .B2(_0238_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_2 _0581_ (.A(_0172_),
    .X(_0239_));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(\updateable_area[24] ),
    .Y(_0240_));
 sky130_fd_sc_hd__clkbuf_4 _0583_ (.A(_0209_),
    .X(_0241_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(net113),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _0585_ (.A(\disruptive_area[24] ),
    .Y(_0243_));
 sky130_fd_sc_hd__or2b_1 _0586_ (.A(_0196_),
    .B_N(\fault_address[24] ),
    .X(_0244_));
 sky130_fd_sc_hd__o221a_1 _0587_ (.A1(_0242_),
    .A2(_0191_),
    .B1(_0243_),
    .B2(_0181_),
    .C1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__o211ai_2 _0588_ (.A1(_0240_),
    .A2(_0241_),
    .B1(_0186_),
    .C1(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__a22o_1 _0589_ (.A1(_0239_),
    .A2(net145),
    .B1(_0231_),
    .B2(_0246_),
    .X(_0163_));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(\disruptive_area[23] ),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(net112),
    .Y(_0248_));
 sky130_fd_sc_hd__buf_4 _0592_ (.A(_0191_),
    .X(_0249_));
 sky130_fd_sc_hd__inv_2 _0593_ (.A(\fault_address[23] ),
    .Y(_0250_));
 sky130_fd_sc_hd__clkbuf_2 _0594_ (.A(_0206_),
    .X(_0251_));
 sky130_fd_sc_hd__inv_2 _0595_ (.A(\updateable_area[23] ),
    .Y(_0252_));
 sky130_fd_sc_hd__o22a_1 _0596_ (.A1(_0250_),
    .A2(_0251_),
    .B1(_0252_),
    .B2(_0216_),
    .X(_0253_));
 sky130_fd_sc_hd__o221ai_4 _0597_ (.A1(_0247_),
    .A2(_0233_),
    .B1(_0248_),
    .B2(_0249_),
    .C1(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__a22o_1 _0598_ (.A1(_0239_),
    .A2(net144),
    .B1(_0231_),
    .B2(_0254_),
    .X(_0162_));
 sky130_fd_sc_hd__inv_2 _0599_ (.A(\updateable_area[22] ),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(net111),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\disruptive_area[22] ),
    .Y(_0257_));
 sky130_fd_sc_hd__or2b_1 _0602_ (.A(_0196_),
    .B_N(\fault_address[22] ),
    .X(_0258_));
 sky130_fd_sc_hd__o221a_1 _0603_ (.A1(_0256_),
    .A2(_0191_),
    .B1(_0257_),
    .B2(_0181_),
    .C1(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__o211ai_4 _0604_ (.A1(_0255_),
    .A2(_0241_),
    .B1(_0186_),
    .C1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__a22o_1 _0605_ (.A1(_0239_),
    .A2(net143),
    .B1(_0231_),
    .B2(_0260_),
    .X(_0161_));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(\disruptive_area[21] ),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _0607_ (.A(net110),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _0608_ (.A(\fault_address[21] ),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _0609_ (.A(\updateable_area[21] ),
    .Y(_0264_));
 sky130_fd_sc_hd__clkbuf_2 _0610_ (.A(_0193_),
    .X(_0265_));
 sky130_fd_sc_hd__o22a_1 _0611_ (.A1(_0263_),
    .A2(_0251_),
    .B1(_0264_),
    .B2(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__o221ai_4 _0612_ (.A1(_0261_),
    .A2(_0233_),
    .B1(_0262_),
    .B2(_0249_),
    .C1(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__a22o_1 _0613_ (.A1(_0239_),
    .A2(net142),
    .B1(_0231_),
    .B2(_0267_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_2 _0614_ (.A(_0174_),
    .X(_0268_));
 sky130_fd_sc_hd__inv_2 _0615_ (.A(\updateable_area[20] ),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _0616_ (.A(net109),
    .Y(_0270_));
 sky130_fd_sc_hd__clkbuf_2 _0617_ (.A(_0190_),
    .X(_0271_));
 sky130_fd_sc_hd__inv_2 _0618_ (.A(\disruptive_area[20] ),
    .Y(_0272_));
 sky130_fd_sc_hd__clkbuf_2 _0619_ (.A(_0179_),
    .X(_0273_));
 sky130_fd_sc_hd__buf_1 _0620_ (.A(_0195_),
    .X(_0274_));
 sky130_fd_sc_hd__or2b_1 _0621_ (.A(_0274_),
    .B_N(\fault_address[20] ),
    .X(_0275_));
 sky130_fd_sc_hd__o221a_1 _0622_ (.A1(_0270_),
    .A2(_0271_),
    .B1(_0272_),
    .B2(_0273_),
    .C1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__o211ai_4 _0623_ (.A1(_0269_),
    .A2(_0241_),
    .B1(_0186_),
    .C1(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__a22o_1 _0624_ (.A1(_0239_),
    .A2(net141),
    .B1(_0268_),
    .B2(_0277_),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_2 _0625_ (.A(_0172_),
    .X(_0278_));
 sky130_fd_sc_hd__inv_2 _0626_ (.A(\disruptive_area[19] ),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _0627_ (.A(net107),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _0628_ (.A(\fault_address[19] ),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0629_ (.A(\updateable_area[19] ),
    .Y(_0282_));
 sky130_fd_sc_hd__o22a_1 _0630_ (.A1(_0281_),
    .A2(_0251_),
    .B1(_0282_),
    .B2(_0265_),
    .X(_0283_));
 sky130_fd_sc_hd__o221ai_4 _0631_ (.A1(_0279_),
    .A2(_0233_),
    .B1(_0280_),
    .B2(_0249_),
    .C1(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__a22o_1 _0632_ (.A1(_0278_),
    .A2(net139),
    .B1(_0268_),
    .B2(_0284_),
    .X(_0158_));
 sky130_fd_sc_hd__inv_2 _0633_ (.A(\updateable_area[18] ),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0634_ (.A(net106),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(\disruptive_area[18] ),
    .Y(_0287_));
 sky130_fd_sc_hd__or2b_1 _0636_ (.A(_0274_),
    .B_N(\fault_address[18] ),
    .X(_0288_));
 sky130_fd_sc_hd__o221a_1 _0637_ (.A1(_0286_),
    .A2(_0271_),
    .B1(_0287_),
    .B2(_0273_),
    .C1(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__o211ai_2 _0638_ (.A1(_0285_),
    .A2(_0241_),
    .B1(_0186_),
    .C1(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__a22o_1 _0639_ (.A1(_0278_),
    .A2(net138),
    .B1(_0268_),
    .B2(_0290_),
    .X(_0157_));
 sky130_fd_sc_hd__inv_2 _0640_ (.A(\updateable_area[17] ),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(net105),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _0642_ (.A(\disruptive_area[17] ),
    .Y(_0293_));
 sky130_fd_sc_hd__or2b_1 _0643_ (.A(_0274_),
    .B_N(\fault_address[17] ),
    .X(_0294_));
 sky130_fd_sc_hd__o221a_1 _0644_ (.A1(_0292_),
    .A2(_0271_),
    .B1(_0293_),
    .B2(_0273_),
    .C1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__o211ai_1 _0645_ (.A1(_0291_),
    .A2(_0241_),
    .B1(_0185_),
    .C1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__a22o_1 _0646_ (.A1(_0278_),
    .A2(net137),
    .B1(_0268_),
    .B2(_0296_),
    .X(_0156_));
 sky130_fd_sc_hd__inv_2 _0647_ (.A(\disruptive_area[16] ),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _0648_ (.A(net104),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _0649_ (.A(\fault_address[16] ),
    .Y(_0299_));
 sky130_fd_sc_hd__inv_2 _0650_ (.A(\updateable_area[16] ),
    .Y(_0300_));
 sky130_fd_sc_hd__o22a_1 _0651_ (.A1(_0299_),
    .A2(_0251_),
    .B1(_0300_),
    .B2(_0265_),
    .X(_0301_));
 sky130_fd_sc_hd__o221ai_2 _0652_ (.A1(_0297_),
    .A2(_0233_),
    .B1(_0298_),
    .B2(_0249_),
    .C1(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__a22o_1 _0653_ (.A1(_0278_),
    .A2(net136),
    .B1(_0268_),
    .B2(_0302_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_2 _0654_ (.A(_0173_),
    .X(_0303_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\disruptive_area[15] ),
    .Y(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _0656_ (.A(_0180_),
    .X(_0305_));
 sky130_fd_sc_hd__inv_2 _0657_ (.A(net103),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _0658_ (.A(\fault_address[15] ),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(\updateable_area[15] ),
    .Y(_0308_));
 sky130_fd_sc_hd__o22a_1 _0660_ (.A1(_0307_),
    .A2(_0251_),
    .B1(_0308_),
    .B2(_0265_),
    .X(_0309_));
 sky130_fd_sc_hd__o221ai_2 _0661_ (.A1(_0304_),
    .A2(_0305_),
    .B1(_0306_),
    .B2(_0249_),
    .C1(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__a22o_1 _0662_ (.A1(_0278_),
    .A2(net135),
    .B1(_0303_),
    .B2(_0310_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_2 _0663_ (.A(_0171_),
    .X(_0311_));
 sky130_fd_sc_hd__inv_2 _0664_ (.A(\disruptive_area[14] ),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(net102),
    .Y(_0313_));
 sky130_fd_sc_hd__clkbuf_4 _0666_ (.A(_0191_),
    .X(_0314_));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(\fault_address[14] ),
    .Y(_0315_));
 sky130_fd_sc_hd__clkbuf_2 _0668_ (.A(_0206_),
    .X(_0316_));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(\updateable_area[14] ),
    .Y(_0317_));
 sky130_fd_sc_hd__o22a_1 _0670_ (.A1(_0315_),
    .A2(_0316_),
    .B1(_0317_),
    .B2(_0265_),
    .X(_0318_));
 sky130_fd_sc_hd__o221ai_2 _0671_ (.A1(_0312_),
    .A2(_0305_),
    .B1(_0313_),
    .B2(_0314_),
    .C1(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__a22o_1 _0672_ (.A1(_0311_),
    .A2(net134),
    .B1(_0303_),
    .B2(_0319_),
    .X(_0153_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(\disruptive_area[13] ),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(net101),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(\fault_address[13] ),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(\updateable_area[13] ),
    .Y(_0323_));
 sky130_fd_sc_hd__clkbuf_2 _0677_ (.A(_0193_),
    .X(_0324_));
 sky130_fd_sc_hd__o22a_1 _0678_ (.A1(_0322_),
    .A2(_0316_),
    .B1(_0323_),
    .B2(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__o221ai_1 _0679_ (.A1(_0320_),
    .A2(_0305_),
    .B1(_0321_),
    .B2(_0314_),
    .C1(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__a22o_1 _0680_ (.A1(_0311_),
    .A2(net133),
    .B1(_0303_),
    .B2(_0326_),
    .X(_0152_));
 sky130_fd_sc_hd__inv_2 _0681_ (.A(\disruptive_area[12] ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(net100),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(\fault_address[12] ),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(\updateable_area[12] ),
    .Y(_0330_));
 sky130_fd_sc_hd__o22a_1 _0685_ (.A1(_0329_),
    .A2(_0316_),
    .B1(_0330_),
    .B2(_0324_),
    .X(_0331_));
 sky130_fd_sc_hd__o221ai_2 _0686_ (.A1(_0327_),
    .A2(_0305_),
    .B1(_0328_),
    .B2(_0314_),
    .C1(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a22o_1 _0687_ (.A1(_0311_),
    .A2(net132),
    .B1(_0303_),
    .B2(_0332_),
    .X(_0151_));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(\disruptive_area[11] ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(net99),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(\fault_address[11] ),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(\updateable_area[11] ),
    .Y(_0336_));
 sky130_fd_sc_hd__o22a_1 _0692_ (.A1(_0335_),
    .A2(_0316_),
    .B1(_0336_),
    .B2(_0324_),
    .X(_0337_));
 sky130_fd_sc_hd__o221ai_4 _0693_ (.A1(_0333_),
    .A2(_0305_),
    .B1(_0334_),
    .B2(_0314_),
    .C1(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__a22o_1 _0694_ (.A1(_0311_),
    .A2(net131),
    .B1(_0303_),
    .B2(_0338_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_2 _0695_ (.A(_0173_),
    .X(_0339_));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(\disruptive_area[10] ),
    .Y(_0340_));
 sky130_fd_sc_hd__clkbuf_4 _0697_ (.A(_0180_),
    .X(_0341_));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(net98),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(\fault_address[10] ),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(\updateable_area[10] ),
    .Y(_0344_));
 sky130_fd_sc_hd__o22a_1 _0701_ (.A1(_0343_),
    .A2(_0316_),
    .B1(_0344_),
    .B2(_0324_),
    .X(_0345_));
 sky130_fd_sc_hd__o221ai_2 _0702_ (.A1(_0340_),
    .A2(_0341_),
    .B1(_0342_),
    .B2(_0314_),
    .C1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a22o_1 _0703_ (.A1(_0311_),
    .A2(net130),
    .B1(_0339_),
    .B2(_0346_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_2 _0704_ (.A(_0171_),
    .X(_0347_));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(\updateable_area[9] ),
    .Y(_0348_));
 sky130_fd_sc_hd__clkbuf_4 _0706_ (.A(_0194_),
    .X(_0349_));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(net128),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(\disruptive_area[9] ),
    .Y(_0351_));
 sky130_fd_sc_hd__or2b_1 _0709_ (.A(_0274_),
    .B_N(\fault_address[9] ),
    .X(_0352_));
 sky130_fd_sc_hd__o221a_1 _0710_ (.A1(_0350_),
    .A2(_0271_),
    .B1(_0351_),
    .B2(_0273_),
    .C1(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__o211ai_2 _0711_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0185_),
    .C1(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__a22o_1 _0712_ (.A1(_0347_),
    .A2(net160),
    .B1(_0339_),
    .B2(_0354_),
    .X(_0148_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(\updateable_area[8] ),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(net127),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(\disruptive_area[8] ),
    .Y(_0357_));
 sky130_fd_sc_hd__or2b_1 _0716_ (.A(_0274_),
    .B_N(\fault_address[8] ),
    .X(_0358_));
 sky130_fd_sc_hd__o221a_1 _0717_ (.A1(_0356_),
    .A2(_0271_),
    .B1(_0357_),
    .B2(_0273_),
    .C1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__o211ai_2 _0718_ (.A1(_0355_),
    .A2(_0349_),
    .B1(_0185_),
    .C1(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__a22o_1 _0719_ (.A1(_0347_),
    .A2(net159),
    .B1(_0339_),
    .B2(_0360_),
    .X(_0147_));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(\disruptive_area[7] ),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(\updateable_area[7] ),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(net126),
    .Y(_0363_));
 sky130_fd_sc_hd__buf_2 _0723_ (.A(_0190_),
    .X(_0364_));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(\fault_address[7] ),
    .Y(_0365_));
 sky130_fd_sc_hd__buf_2 _0725_ (.A(_0195_),
    .X(_0366_));
 sky130_fd_sc_hd__or4_4 _0726_ (.A(net8),
    .B(_0177_),
    .C(_0183_),
    .D(_0188_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_2 _0727_ (.A(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__or2b_1 _0728_ (.A(_0368_),
    .B_N(\fault_status[7] ),
    .X(_0369_));
 sky130_fd_sc_hd__o221a_1 _0729_ (.A1(_0363_),
    .A2(_0364_),
    .B1(_0365_),
    .B2(_0366_),
    .C1(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__o221ai_2 _0730_ (.A1(_0361_),
    .A2(_0341_),
    .B1(_0362_),
    .B2(_0349_),
    .C1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(_0347_),
    .A2(net158),
    .B1(_0339_),
    .B2(_0371_),
    .X(_0146_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(\disruptive_area[6] ),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(\updateable_area[6] ),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(net125),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(\fault_address[6] ),
    .Y(_0375_));
 sky130_fd_sc_hd__or2b_1 _0736_ (.A(_0368_),
    .B_N(\fault_status[6] ),
    .X(_0376_));
 sky130_fd_sc_hd__o221a_1 _0737_ (.A1(_0374_),
    .A2(_0364_),
    .B1(_0375_),
    .B2(_0366_),
    .C1(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__o221ai_2 _0738_ (.A1(_0372_),
    .A2(_0341_),
    .B1(_0373_),
    .B2(_0349_),
    .C1(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(_0347_),
    .A2(net157),
    .B1(_0339_),
    .B2(_0378_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_2 _0740_ (.A(_0173_),
    .X(_0379_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(\disruptive_area[5] ),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(\updateable_area[5] ),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(net124),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(\fault_address[5] ),
    .Y(_0383_));
 sky130_fd_sc_hd__or2b_1 _0745_ (.A(_0367_),
    .B_N(\fault_status[5] ),
    .X(_0384_));
 sky130_fd_sc_hd__o221a_1 _0746_ (.A1(_0382_),
    .A2(_0364_),
    .B1(_0383_),
    .B2(_0366_),
    .C1(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__o221ai_2 _0747_ (.A1(_0380_),
    .A2(_0341_),
    .B1(_0381_),
    .B2(_0349_),
    .C1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a22o_1 _0748_ (.A1(_0347_),
    .A2(net156),
    .B1(_0379_),
    .B2(_0386_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_2 _0749_ (.A(_0171_),
    .X(_0387_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(\disruptive_area[4] ),
    .Y(_0388_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(\updateable_area[4] ),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(net123),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(\fault_address[4] ),
    .Y(_0391_));
 sky130_fd_sc_hd__or2b_1 _0754_ (.A(_0367_),
    .B_N(\fault_status[4] ),
    .X(_0392_));
 sky130_fd_sc_hd__o221a_1 _0755_ (.A1(_0390_),
    .A2(_0364_),
    .B1(_0391_),
    .B2(_0366_),
    .C1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__o221ai_2 _0756_ (.A1(_0388_),
    .A2(_0341_),
    .B1(_0389_),
    .B2(_0209_),
    .C1(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a22o_1 _0757_ (.A1(_0387_),
    .A2(net155),
    .B1(_0379_),
    .B2(_0394_),
    .X(_0143_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(\disruptive_area[3] ),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(\updateable_area[3] ),
    .Y(_0396_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(net122),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(\fault_address[3] ),
    .Y(_0398_));
 sky130_fd_sc_hd__or2b_1 _0762_ (.A(_0367_),
    .B_N(\fault_status[3] ),
    .X(_0399_));
 sky130_fd_sc_hd__o221a_1 _0763_ (.A1(_0397_),
    .A2(_0364_),
    .B1(_0398_),
    .B2(_0196_),
    .C1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__o221ai_2 _0764_ (.A1(_0395_),
    .A2(_0181_),
    .B1(_0396_),
    .B2(_0209_),
    .C1(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a22o_1 _0765_ (.A1(_0387_),
    .A2(net154),
    .B1(_0379_),
    .B2(_0401_),
    .X(_0142_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(\fault_status[2] ),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(net119),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(\updateable_area[2] ),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(\cache_control[2] ),
    .Y(_0405_));
 sky130_fd_sc_hd__or3_4 _0770_ (.A(_0183_),
    .B(_0189_),
    .C(_0184_),
    .X(_0406_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(\fault_address[2] ),
    .Y(_0407_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(\disruptive_area[2] ),
    .Y(_0408_));
 sky130_fd_sc_hd__o22a_1 _0773_ (.A1(_0407_),
    .A2(_0206_),
    .B1(_0408_),
    .B2(_0180_),
    .X(_0409_));
 sky130_fd_sc_hd__o221a_1 _0774_ (.A1(_0404_),
    .A2(_0194_),
    .B1(_0405_),
    .B2(_0406_),
    .C1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__o221ai_2 _0775_ (.A1(_0402_),
    .A2(_0368_),
    .B1(_0403_),
    .B2(_0203_),
    .C1(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__a22o_1 _0776_ (.A1(_0387_),
    .A2(net151),
    .B1(_0379_),
    .B2(_0411_),
    .X(_0141_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(\fault_status[1] ),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(net108),
    .Y(_0413_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(\updateable_area[1] ),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(\cache_control[1] ),
    .Y(_0415_));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(\fault_address[1] ),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(\disruptive_area[1] ),
    .Y(_0417_));
 sky130_fd_sc_hd__o22a_1 _0783_ (.A1(_0416_),
    .A2(_0206_),
    .B1(_0417_),
    .B2(_0179_),
    .X(_0418_));
 sky130_fd_sc_hd__o221a_1 _0784_ (.A1(_0414_),
    .A2(_0194_),
    .B1(_0415_),
    .B2(_0406_),
    .C1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__o221ai_2 _0785_ (.A1(_0412_),
    .A2(_0368_),
    .B1(_0413_),
    .B2(_0203_),
    .C1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__a22o_1 _0786_ (.A1(_0387_),
    .A2(net140),
    .B1(_0379_),
    .B2(_0420_),
    .X(_0140_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(net97),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(\updateable_area[0] ),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(\fault_address[0] ),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(net95),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(\fault_status[0] ),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(\disruptive_area[0] ),
    .Y(_0426_));
 sky130_fd_sc_hd__o22a_1 _0793_ (.A1(_0425_),
    .A2(_0368_),
    .B1(_0426_),
    .B2(_0179_),
    .X(_0427_));
 sky130_fd_sc_hd__o221a_1 _0794_ (.A1(_0423_),
    .A2(_0196_),
    .B1(_0424_),
    .B2(_0406_),
    .C1(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__o221ai_1 _0795_ (.A1(_0421_),
    .A2(_0203_),
    .B1(_0422_),
    .B2(_0209_),
    .C1(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__a22o_1 _0796_ (.A1(_0387_),
    .A2(net129),
    .B1(_0174_),
    .B2(_0429_),
    .X(_0139_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(net20),
    .Y(_0430_));
 sky130_fd_sc_hd__or4_4 _0798_ (.A(_0171_),
    .B(net19),
    .C(_0430_),
    .D(_0179_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_2 _0799_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_2 _0800_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(_0431_),
    .Y(_0434_));
 sky130_fd_sc_hd__clkbuf_2 _0802_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_2 _0803_ (.A(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(\disruptive_area[31] ),
    .A2(_0433_),
    .B1(net45),
    .B2(_0436_),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(\disruptive_area[30] ),
    .A2(_0433_),
    .B1(net44),
    .B2(_0436_),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _0806_ (.A1(\disruptive_area[29] ),
    .A2(_0433_),
    .B1(net42),
    .B2(_0436_),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _0807_ (.A1(\disruptive_area[28] ),
    .A2(_0433_),
    .B1(net41),
    .B2(_0436_),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(\disruptive_area[27] ),
    .A2(_0433_),
    .B1(net40),
    .B2(_0436_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_2 _0809_ (.A(_0432_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_2 _0810_ (.A(_0435_),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _0811_ (.A1(\disruptive_area[26] ),
    .A2(_0437_),
    .B1(net39),
    .B2(_0438_),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0812_ (.A1(\disruptive_area[25] ),
    .A2(_0437_),
    .B1(net38),
    .B2(_0438_),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _0813_ (.A1(\disruptive_area[24] ),
    .A2(_0437_),
    .B1(net37),
    .B2(_0438_),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(\disruptive_area[23] ),
    .A2(_0437_),
    .B1(net36),
    .B2(_0438_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _0815_ (.A1(\disruptive_area[22] ),
    .A2(_0437_),
    .B1(net35),
    .B2(_0438_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_2 _0816_ (.A(_0432_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_2 _0817_ (.A(_0435_),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _0818_ (.A1(\disruptive_area[21] ),
    .A2(_0439_),
    .B1(net34),
    .B2(_0440_),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _0819_ (.A1(\disruptive_area[20] ),
    .A2(_0439_),
    .B1(net33),
    .B2(_0440_),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _0820_ (.A1(\disruptive_area[19] ),
    .A2(_0439_),
    .B1(net31),
    .B2(_0440_),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _0821_ (.A1(\disruptive_area[18] ),
    .A2(_0439_),
    .B1(net30),
    .B2(_0440_),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(\disruptive_area[17] ),
    .A2(_0439_),
    .B1(net29),
    .B2(_0440_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_2 _0823_ (.A(_0431_),
    .X(_0441_));
 sky130_fd_sc_hd__buf_1 _0824_ (.A(_0434_),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_1 _0825_ (.A1(\disruptive_area[16] ),
    .A2(_0441_),
    .B1(net28),
    .B2(_0442_),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(\disruptive_area[15] ),
    .A2(_0441_),
    .B1(net27),
    .B2(_0442_),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _0827_ (.A1(\disruptive_area[14] ),
    .A2(_0441_),
    .B1(net26),
    .B2(_0442_),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(\disruptive_area[13] ),
    .A2(_0441_),
    .B1(net25),
    .B2(_0442_),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _0829_ (.A1(\disruptive_area[12] ),
    .A2(_0441_),
    .B1(net24),
    .B2(_0442_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_2 _0830_ (.A(_0431_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_2 _0831_ (.A(_0434_),
    .X(_0444_));
 sky130_fd_sc_hd__a22o_1 _0832_ (.A1(\disruptive_area[11] ),
    .A2(_0443_),
    .B1(net23),
    .B2(_0444_),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(\disruptive_area[10] ),
    .A2(_0443_),
    .B1(net22),
    .B2(_0444_),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _0834_ (.A1(\disruptive_area[9] ),
    .A2(_0443_),
    .B1(net52),
    .B2(_0444_),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_1 _0835_ (.A1(\disruptive_area[8] ),
    .A2(_0443_),
    .B1(net51),
    .B2(_0444_),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _0836_ (.A1(\disruptive_area[7] ),
    .A2(_0443_),
    .B1(net50),
    .B2(_0444_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_2 _0837_ (.A(_0431_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_2 _0838_ (.A(_0434_),
    .X(_0446_));
 sky130_fd_sc_hd__a22o_1 _0839_ (.A1(\disruptive_area[6] ),
    .A2(_0445_),
    .B1(net49),
    .B2(_0446_),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _0840_ (.A1(\disruptive_area[5] ),
    .A2(_0445_),
    .B1(net48),
    .B2(_0446_),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(\disruptive_area[4] ),
    .A2(_0445_),
    .B1(net47),
    .B2(_0446_),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _0842_ (.A1(\disruptive_area[3] ),
    .A2(_0445_),
    .B1(net46),
    .B2(_0446_),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _0843_ (.A1(\disruptive_area[2] ),
    .A2(_0445_),
    .B1(net43),
    .B2(_0446_),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _0844_ (.A1(\disruptive_area[1] ),
    .A2(_0432_),
    .B1(net32),
    .B2(_0435_),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _0845_ (.A1(\disruptive_area[0] ),
    .A2(_0432_),
    .B1(net21),
    .B2(_0435_),
    .X(_0107_));
 sky130_fd_sc_hd__or4_4 _0846_ (.A(net53),
    .B(net19),
    .C(_0430_),
    .D(_0193_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_2 _0847_ (.A(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_2 _0848_ (.A(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__inv_2 _0849_ (.A(_0447_),
    .Y(_0450_));
 sky130_fd_sc_hd__clkbuf_2 _0850_ (.A(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_2 _0851_ (.A(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(\updateable_area[31] ),
    .A2(_0449_),
    .B1(net45),
    .B2(_0452_),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_1 _0853_ (.A1(\updateable_area[30] ),
    .A2(_0449_),
    .B1(net44),
    .B2(_0452_),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(\updateable_area[29] ),
    .A2(_0449_),
    .B1(net42),
    .B2(_0452_),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_1 _0855_ (.A1(\updateable_area[28] ),
    .A2(_0449_),
    .B1(net41),
    .B2(_0452_),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(\updateable_area[27] ),
    .A2(_0449_),
    .B1(net40),
    .B2(_0452_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_2 _0857_ (.A(_0448_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_2 _0858_ (.A(_0451_),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(\updateable_area[26] ),
    .A2(_0453_),
    .B1(net39),
    .B2(_0454_),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_1 _0860_ (.A1(\updateable_area[25] ),
    .A2(_0453_),
    .B1(net38),
    .B2(_0454_),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _0861_ (.A1(\updateable_area[24] ),
    .A2(_0453_),
    .B1(net37),
    .B2(_0454_),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _0862_ (.A1(\updateable_area[23] ),
    .A2(_0453_),
    .B1(net36),
    .B2(_0454_),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_1 _0863_ (.A1(\updateable_area[22] ),
    .A2(_0453_),
    .B1(net35),
    .B2(_0454_),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_2 _0864_ (.A(_0448_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_2 _0865_ (.A(_0451_),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _0866_ (.A1(\updateable_area[21] ),
    .A2(_0455_),
    .B1(net34),
    .B2(_0456_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _0867_ (.A1(\updateable_area[20] ),
    .A2(_0455_),
    .B1(net33),
    .B2(_0456_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _0868_ (.A1(\updateable_area[19] ),
    .A2(_0455_),
    .B1(net31),
    .B2(_0456_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _0869_ (.A1(\updateable_area[18] ),
    .A2(_0455_),
    .B1(net30),
    .B2(_0456_),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_1 _0870_ (.A1(\updateable_area[17] ),
    .A2(_0455_),
    .B1(net29),
    .B2(_0456_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_2 _0871_ (.A(_0447_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_2 _0872_ (.A(_0450_),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _0873_ (.A1(\updateable_area[16] ),
    .A2(_0457_),
    .B1(net28),
    .B2(_0458_),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _0874_ (.A1(\updateable_area[15] ),
    .A2(_0457_),
    .B1(net27),
    .B2(_0458_),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _0875_ (.A1(\updateable_area[14] ),
    .A2(_0457_),
    .B1(net26),
    .B2(_0458_),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _0876_ (.A1(\updateable_area[13] ),
    .A2(_0457_),
    .B1(net25),
    .B2(_0458_),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _0877_ (.A1(\updateable_area[12] ),
    .A2(_0457_),
    .B1(net24),
    .B2(_0458_),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_2 _0878_ (.A(_0447_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_2 _0879_ (.A(_0450_),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _0880_ (.A1(\updateable_area[11] ),
    .A2(_0459_),
    .B1(net23),
    .B2(_0460_),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _0881_ (.A1(\updateable_area[10] ),
    .A2(_0459_),
    .B1(net22),
    .B2(_0460_),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _0882_ (.A1(\updateable_area[9] ),
    .A2(_0459_),
    .B1(net52),
    .B2(_0460_),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _0883_ (.A1(\updateable_area[8] ),
    .A2(_0459_),
    .B1(net51),
    .B2(_0460_),
    .X(_0083_));
 sky130_fd_sc_hd__a22o_1 _0884_ (.A1(\updateable_area[7] ),
    .A2(_0459_),
    .B1(net50),
    .B2(_0460_),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_2 _0885_ (.A(_0447_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_2 _0886_ (.A(_0450_),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _0887_ (.A1(\updateable_area[6] ),
    .A2(_0461_),
    .B1(net49),
    .B2(_0462_),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_1 _0888_ (.A1(\updateable_area[5] ),
    .A2(_0461_),
    .B1(net48),
    .B2(_0462_),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _0889_ (.A1(\updateable_area[4] ),
    .A2(_0461_),
    .B1(net47),
    .B2(_0462_),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _0890_ (.A1(\updateable_area[3] ),
    .A2(_0461_),
    .B1(net46),
    .B2(_0462_),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _0891_ (.A1(\updateable_area[2] ),
    .A2(_0461_),
    .B1(net43),
    .B2(_0462_),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _0892_ (.A1(\updateable_area[1] ),
    .A2(_0448_),
    .B1(net32),
    .B2(_0451_),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_1 _0893_ (.A1(\updateable_area[0] ),
    .A2(_0448_),
    .B1(net21),
    .B2(_0451_),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_2 _0894_ (.A(_0173_),
    .B(net54),
    .Y(_0463_));
 sky130_fd_sc_hd__buf_2 _0895_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_2 _0896_ (.A(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__inv_2 _0897_ (.A(_0463_),
    .Y(_0466_));
 sky130_fd_sc_hd__buf_2 _0898_ (.A(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_2 _0899_ (.A(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _0900_ (.A1(\fault_address[31] ),
    .A2(_0465_),
    .B1(net79),
    .B2(_0468_),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_1 _0901_ (.A1(\fault_address[30] ),
    .A2(_0465_),
    .B1(net78),
    .B2(_0468_),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _0902_ (.A1(\fault_address[29] ),
    .A2(_0465_),
    .B1(net76),
    .B2(_0468_),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_1 _0903_ (.A1(\fault_address[28] ),
    .A2(_0465_),
    .B1(net75),
    .B2(_0468_),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _0904_ (.A1(\fault_address[27] ),
    .A2(_0465_),
    .B1(net74),
    .B2(_0468_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_2 _0905_ (.A(_0464_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_2 _0906_ (.A(_0467_),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _0907_ (.A1(\fault_address[26] ),
    .A2(_0469_),
    .B1(net73),
    .B2(_0470_),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _0908_ (.A1(\fault_address[25] ),
    .A2(_0469_),
    .B1(net72),
    .B2(_0470_),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _0909_ (.A1(\fault_address[24] ),
    .A2(_0469_),
    .B1(net71),
    .B2(_0470_),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _0910_ (.A1(\fault_address[23] ),
    .A2(_0469_),
    .B1(net70),
    .B2(_0470_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _0911_ (.A1(\fault_address[22] ),
    .A2(_0469_),
    .B1(net69),
    .B2(_0470_),
    .X(_0065_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0912_ (.A(_0464_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_2 _0913_ (.A(_0467_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(\fault_address[21] ),
    .A2(_0471_),
    .B1(net68),
    .B2(_0472_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _0915_ (.A1(\fault_address[20] ),
    .A2(_0471_),
    .B1(net67),
    .B2(_0472_),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _0916_ (.A1(\fault_address[19] ),
    .A2(_0471_),
    .B1(net65),
    .B2(_0472_),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _0917_ (.A1(\fault_address[18] ),
    .A2(_0471_),
    .B1(net64),
    .B2(_0472_),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_1 _0918_ (.A1(\fault_address[17] ),
    .A2(_0471_),
    .B1(net63),
    .B2(_0472_),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_2 _0919_ (.A(_0464_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_2 _0920_ (.A(_0467_),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _0921_ (.A1(\fault_address[16] ),
    .A2(_0473_),
    .B1(net62),
    .B2(_0474_),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _0922_ (.A1(\fault_address[15] ),
    .A2(_0473_),
    .B1(net61),
    .B2(_0474_),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _0923_ (.A1(\fault_address[14] ),
    .A2(_0473_),
    .B1(net60),
    .B2(_0474_),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_1 _0924_ (.A1(\fault_address[13] ),
    .A2(_0473_),
    .B1(net59),
    .B2(_0474_),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _0925_ (.A1(\fault_address[12] ),
    .A2(_0473_),
    .B1(net58),
    .B2(_0474_),
    .X(_0055_));
 sky130_fd_sc_hd__clkbuf_2 _0926_ (.A(_0464_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_2 _0927_ (.A(_0467_),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _0928_ (.A1(\fault_address[11] ),
    .A2(_0475_),
    .B1(net57),
    .B2(_0476_),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _0929_ (.A1(\fault_address[10] ),
    .A2(_0475_),
    .B1(net56),
    .B2(_0476_),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _0930_ (.A1(\fault_address[9] ),
    .A2(_0475_),
    .B1(net86),
    .B2(_0476_),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _0931_ (.A1(\fault_address[8] ),
    .A2(_0475_),
    .B1(net85),
    .B2(_0476_),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _0932_ (.A1(\fault_address[7] ),
    .A2(_0475_),
    .B1(net84),
    .B2(_0476_),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_2 _0933_ (.A(_0463_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_2 _0934_ (.A(_0466_),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _0935_ (.A1(\fault_address[6] ),
    .A2(_0477_),
    .B1(net83),
    .B2(_0478_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _0936_ (.A1(\fault_address[5] ),
    .A2(_0477_),
    .B1(net82),
    .B2(_0478_),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _0937_ (.A1(\fault_address[4] ),
    .A2(_0477_),
    .B1(net81),
    .B2(_0478_),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _0938_ (.A1(\fault_address[3] ),
    .A2(_0477_),
    .B1(net80),
    .B2(_0478_),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_1 _0939_ (.A1(\fault_address[2] ),
    .A2(_0477_),
    .B1(net77),
    .B2(_0478_),
    .X(_0045_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0940_ (.A(_0463_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_2 _0941_ (.A(_0466_),
    .X(_0480_));
 sky130_fd_sc_hd__a22o_1 _0942_ (.A1(\fault_address[1] ),
    .A2(_0479_),
    .B1(net66),
    .B2(_0480_),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_1 _0943_ (.A1(\fault_address[0] ),
    .A2(_0479_),
    .B1(net55),
    .B2(_0480_),
    .X(_0043_));
 sky130_fd_sc_hd__or4_4 _0944_ (.A(net53),
    .B(net19),
    .C(_0430_),
    .D(_0184_),
    .X(_0481_));
 sky130_fd_sc_hd__or3_4 _0945_ (.A(_0178_),
    .B(_0189_),
    .C(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_2 _0946_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_2 _0947_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(_0482_),
    .Y(_0485_));
 sky130_fd_sc_hd__clkbuf_2 _0949_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_2 _0950_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _0951_ (.A1(net121),
    .A2(_0484_),
    .B1(net45),
    .B2(_0487_),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _0952_ (.A1(net120),
    .A2(_0484_),
    .B1(net44),
    .B2(_0487_),
    .X(_0041_));
 sky130_fd_sc_hd__a22o_1 _0953_ (.A1(net118),
    .A2(_0484_),
    .B1(net42),
    .B2(_0487_),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _0954_ (.A1(net117),
    .A2(_0484_),
    .B1(net41),
    .B2(_0487_),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _0955_ (.A1(net116),
    .A2(_0484_),
    .B1(net40),
    .B2(_0487_),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_2 _0956_ (.A(_0483_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_2 _0957_ (.A(_0486_),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _0958_ (.A1(net115),
    .A2(_0488_),
    .B1(net39),
    .B2(_0489_),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _0959_ (.A1(net114),
    .A2(_0488_),
    .B1(net38),
    .B2(_0489_),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _0960_ (.A1(net113),
    .A2(_0488_),
    .B1(net37),
    .B2(_0489_),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _0961_ (.A1(net112),
    .A2(_0488_),
    .B1(net36),
    .B2(_0489_),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _0962_ (.A1(net111),
    .A2(_0488_),
    .B1(net35),
    .B2(_0489_),
    .X(_0033_));
 sky130_fd_sc_hd__clkbuf_2 _0963_ (.A(_0483_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_2 _0964_ (.A(_0486_),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _0965_ (.A1(net110),
    .A2(_0490_),
    .B1(net34),
    .B2(_0491_),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _0966_ (.A1(net109),
    .A2(_0490_),
    .B1(net33),
    .B2(_0491_),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _0967_ (.A1(net107),
    .A2(_0490_),
    .B1(net31),
    .B2(_0491_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _0968_ (.A1(net106),
    .A2(_0490_),
    .B1(net30),
    .B2(_0491_),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _0969_ (.A1(net105),
    .A2(_0490_),
    .B1(net29),
    .B2(_0491_),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_2 _0970_ (.A(_0482_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_2 _0971_ (.A(_0485_),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _0972_ (.A1(net104),
    .A2(_0492_),
    .B1(net28),
    .B2(_0493_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_1 _0973_ (.A1(net103),
    .A2(_0492_),
    .B1(net27),
    .B2(_0493_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_1 _0974_ (.A1(net102),
    .A2(_0492_),
    .B1(net26),
    .B2(_0493_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _0975_ (.A1(net101),
    .A2(_0492_),
    .B1(net25),
    .B2(_0493_),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_1 _0976_ (.A1(net100),
    .A2(_0492_),
    .B1(net24),
    .B2(_0493_),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_2 _0977_ (.A(_0482_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_2 _0978_ (.A(_0485_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _0979_ (.A1(net99),
    .A2(_0494_),
    .B1(net23),
    .B2(_0495_),
    .X(_0022_));
 sky130_fd_sc_hd__a22o_1 _0980_ (.A1(net98),
    .A2(_0494_),
    .B1(net22),
    .B2(_0495_),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_1 _0981_ (.A1(net128),
    .A2(_0494_),
    .B1(net52),
    .B2(_0495_),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_1 _0982_ (.A1(net127),
    .A2(_0494_),
    .B1(net51),
    .B2(_0495_),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _0983_ (.A1(net126),
    .A2(_0494_),
    .B1(net50),
    .B2(_0495_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_2 _0984_ (.A(_0482_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_2 _0985_ (.A(_0485_),
    .X(_0497_));
 sky130_fd_sc_hd__a22o_1 _0986_ (.A1(net125),
    .A2(_0496_),
    .B1(net49),
    .B2(_0497_),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _0987_ (.A1(net124),
    .A2(_0496_),
    .B1(net48),
    .B2(_0497_),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _0988_ (.A1(net123),
    .A2(_0496_),
    .B1(net47),
    .B2(_0497_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _0989_ (.A1(net122),
    .A2(_0496_),
    .B1(net46),
    .B2(_0497_),
    .X(_0014_));
 sky130_fd_sc_hd__a22o_1 _0990_ (.A1(net119),
    .A2(_0496_),
    .B1(net43),
    .B2(_0497_),
    .X(_0013_));
 sky130_fd_sc_hd__a22o_1 _0991_ (.A1(net108),
    .A2(_0483_),
    .B1(net32),
    .B2(_0486_),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_1 _0992_ (.A1(net97),
    .A2(_0483_),
    .B1(net21),
    .B2(_0486_),
    .X(_0011_));
 sky130_fd_sc_hd__or3_4 _0993_ (.A(_0183_),
    .B(_0189_),
    .C(_0481_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(net43),
    .A1(\cache_control[2] ),
    .S(_0498_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(net32),
    .A1(\cache_control[1] ),
    .S(_0498_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net21),
    .A1(net95),
    .S(_0498_),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_1 _0997_ (.A1(\fault_status[7] ),
    .A2(_0479_),
    .B1(net94),
    .B2(_0480_),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_1 _0998_ (.A1(\fault_status[6] ),
    .A2(_0479_),
    .B1(net93),
    .B2(_0480_),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _0999_ (.A1(\fault_status[5] ),
    .A2(_0479_),
    .B1(net92),
    .B2(_0480_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_2 _1000_ (.A(_0463_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_2 _1001_ (.A(_0466_),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _1002_ (.A1(\fault_status[4] ),
    .A2(_0499_),
    .B1(net91),
    .B2(_0500_),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _1003_ (.A1(\fault_status[3] ),
    .A2(_0499_),
    .B1(net90),
    .B2(_0500_),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _1004_ (.A1(\fault_status[2] ),
    .A2(_0499_),
    .B1(net89),
    .B2(_0500_),
    .X(_0002_));
 sky130_fd_sc_hd__a22o_1 _1005_ (.A1(\fault_status[1] ),
    .A2(_0499_),
    .B1(net88),
    .B2(_0500_),
    .X(_0001_));
 sky130_fd_sc_hd__a22o_1 _1006_ (.A1(\fault_status[0] ),
    .A2(_0499_),
    .B1(net87),
    .B2(_0500_),
    .X(_0000_));
 sky130_fd_sc_hd__nor3_4 _1007_ (.A(_0178_),
    .B(net6),
    .C(_0481_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(\disruptive_area[31] ),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(net121),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _1010_ (.A(\fault_address[31] ),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(\updateable_area[31] ),
    .Y(_0504_));
 sky130_fd_sc_hd__o22a_1 _1012_ (.A1(_0503_),
    .A2(_0366_),
    .B1(_0504_),
    .B2(_0324_),
    .X(_0505_));
 sky130_fd_sc_hd__o221ai_2 _1013_ (.A1(_0501_),
    .A2(_0181_),
    .B1(_0502_),
    .B2(_0203_),
    .C1(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__a22o_1 _1014_ (.A1(_0172_),
    .A2(net153),
    .B1(_0174_),
    .B2(_0506_),
    .X(_0170_));
 sky130_fd_sc_hd__buf_2 _1015_ (.A(net97),
    .X(\cacheable_area[0] ));
 sky130_fd_sc_hd__buf_2 _1016_ (.A(net108),
    .X(\cacheable_area[1] ));
 sky130_fd_sc_hd__buf_2 _1017_ (.A(net119),
    .X(\cacheable_area[2] ));
 sky130_fd_sc_hd__buf_2 _1018_ (.A(net122),
    .X(\cacheable_area[3] ));
 sky130_fd_sc_hd__buf_2 _1019_ (.A(net123),
    .X(\cacheable_area[4] ));
 sky130_fd_sc_hd__buf_2 _1020_ (.A(net124),
    .X(\cacheable_area[5] ));
 sky130_fd_sc_hd__buf_2 _1021_ (.A(net125),
    .X(\cacheable_area[6] ));
 sky130_fd_sc_hd__buf_2 _1022_ (.A(net126),
    .X(\cacheable_area[7] ));
 sky130_fd_sc_hd__buf_2 _1023_ (.A(net127),
    .X(\cacheable_area[8] ));
 sky130_fd_sc_hd__buf_2 _1024_ (.A(net128),
    .X(\cacheable_area[9] ));
 sky130_fd_sc_hd__buf_2 _1025_ (.A(net98),
    .X(\cacheable_area[10] ));
 sky130_fd_sc_hd__buf_2 _1026_ (.A(net99),
    .X(\cacheable_area[11] ));
 sky130_fd_sc_hd__buf_2 _1027_ (.A(net100),
    .X(\cacheable_area[12] ));
 sky130_fd_sc_hd__buf_2 _1028_ (.A(net101),
    .X(\cacheable_area[13] ));
 sky130_fd_sc_hd__buf_2 _1029_ (.A(net102),
    .X(\cacheable_area[14] ));
 sky130_fd_sc_hd__buf_2 _1030_ (.A(net103),
    .X(\cacheable_area[15] ));
 sky130_fd_sc_hd__buf_2 _1031_ (.A(net104),
    .X(\cacheable_area[16] ));
 sky130_fd_sc_hd__buf_2 _1032_ (.A(net105),
    .X(\cacheable_area[17] ));
 sky130_fd_sc_hd__buf_2 _1033_ (.A(net106),
    .X(\cacheable_area[18] ));
 sky130_fd_sc_hd__buf_2 _1034_ (.A(net107),
    .X(\cacheable_area[19] ));
 sky130_fd_sc_hd__buf_2 _1035_ (.A(net109),
    .X(\cacheable_area[20] ));
 sky130_fd_sc_hd__buf_2 _1036_ (.A(net110),
    .X(\cacheable_area[21] ));
 sky130_fd_sc_hd__buf_2 _1037_ (.A(net111),
    .X(\cacheable_area[22] ));
 sky130_fd_sc_hd__buf_2 _1038_ (.A(net112),
    .X(\cacheable_area[23] ));
 sky130_fd_sc_hd__buf_2 _1039_ (.A(net113),
    .X(\cacheable_area[24] ));
 sky130_fd_sc_hd__buf_2 _1040_ (.A(net114),
    .X(\cacheable_area[25] ));
 sky130_fd_sc_hd__buf_2 _1041_ (.A(net115),
    .X(\cacheable_area[26] ));
 sky130_fd_sc_hd__buf_2 _1042_ (.A(net116),
    .X(\cacheable_area[27] ));
 sky130_fd_sc_hd__buf_2 _1043_ (.A(net117),
    .X(\cacheable_area[28] ));
 sky130_fd_sc_hd__buf_2 _1044_ (.A(net118),
    .X(\cacheable_area[29] ));
 sky130_fd_sc_hd__buf_2 _1045_ (.A(net120),
    .X(\cacheable_area[30] ));
 sky130_fd_sc_hd__buf_2 _1046_ (.A(net121),
    .X(\cacheable_area[31] ));
 sky130_fd_sc_hd__buf_2 _1047_ (.A(net95),
    .X(\cache_control[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.D(_0000_),
    .Q(\fault_status[0] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.D(_0001_),
    .Q(\fault_status[1] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.D(_0002_),
    .Q(\fault_status[2] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.D(_0003_),
    .Q(\fault_status[3] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.D(_0004_),
    .Q(\fault_status[4] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.D(_0005_),
    .Q(\fault_status[5] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.D(_0006_),
    .Q(\fault_status[6] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.D(_0007_),
    .Q(\fault_status[7] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1056_ (.D(_0008_),
    .Q(net95),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.D(_0009_),
    .Q(\cache_control[1] ),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.D(_0010_),
    .Q(\cache_control[2] ),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1059_ (.D(_0011_),
    .Q(net97),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1060_ (.D(_0012_),
    .Q(net108),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1061_ (.D(_0013_),
    .Q(net119),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1062_ (.D(_0014_),
    .Q(net122),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1063_ (.D(_0015_),
    .Q(net123),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1064_ (.D(_0016_),
    .Q(net124),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1065_ (.D(_0017_),
    .Q(net125),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.D(_0018_),
    .Q(net126),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.D(_0019_),
    .Q(net127),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.D(_0020_),
    .Q(net128),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1069_ (.D(_0021_),
    .Q(net98),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.D(_0022_),
    .Q(net99),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1071_ (.D(_0023_),
    .Q(net100),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.D(_0024_),
    .Q(net101),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1073_ (.D(_0025_),
    .Q(net102),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1074_ (.D(_0026_),
    .Q(net103),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.D(_0027_),
    .Q(net104),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.D(_0028_),
    .Q(net105),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1077_ (.D(_0029_),
    .Q(net106),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1078_ (.D(_0030_),
    .Q(net107),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1079_ (.D(_0031_),
    .Q(net109),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.D(_0032_),
    .Q(net110),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1081_ (.D(_0033_),
    .Q(net111),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1082_ (.D(_0034_),
    .Q(net112),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.D(_0035_),
    .Q(net113),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.D(_0036_),
    .Q(net114),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1085_ (.D(_0037_),
    .Q(net115),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.D(_0038_),
    .Q(net116),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1087_ (.D(_0039_),
    .Q(net117),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1088_ (.D(_0040_),
    .Q(net118),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1089_ (.D(_0041_),
    .Q(net120),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1090_ (.D(_0042_),
    .Q(net121),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.D(_0043_),
    .Q(\fault_address[0] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.D(_0044_),
    .Q(\fault_address[1] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.D(_0045_),
    .Q(\fault_address[2] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.D(_0046_),
    .Q(\fault_address[3] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.D(_0047_),
    .Q(\fault_address[4] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.D(_0048_),
    .Q(\fault_address[5] ),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.D(_0049_),
    .Q(\fault_address[6] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.D(_0050_),
    .Q(\fault_address[7] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.D(_0051_),
    .Q(\fault_address[8] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.D(_0052_),
    .Q(\fault_address[9] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.D(_0053_),
    .Q(\fault_address[10] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.D(_0054_),
    .Q(\fault_address[11] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.D(_0055_),
    .Q(\fault_address[12] ),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.D(_0056_),
    .Q(\fault_address[13] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.D(_0057_),
    .Q(\fault_address[14] ),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.D(_0058_),
    .Q(\fault_address[15] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.D(_0059_),
    .Q(\fault_address[16] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.D(_0060_),
    .Q(\fault_address[17] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.D(_0061_),
    .Q(\fault_address[18] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.D(_0062_),
    .Q(\fault_address[19] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.D(_0063_),
    .Q(\fault_address[20] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.D(_0064_),
    .Q(\fault_address[21] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.D(_0065_),
    .Q(\fault_address[22] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.D(_0066_),
    .Q(\fault_address[23] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.D(_0067_),
    .Q(\fault_address[24] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.D(_0068_),
    .Q(\fault_address[25] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.D(_0069_),
    .Q(\fault_address[26] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.D(_0070_),
    .Q(\fault_address[27] ),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.D(_0071_),
    .Q(\fault_address[28] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.D(_0072_),
    .Q(\fault_address[29] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.D(_0073_),
    .Q(\fault_address[30] ),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.D(_0074_),
    .Q(\fault_address[31] ),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.D(_0075_),
    .Q(\updateable_area[0] ),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.D(_0076_),
    .Q(\updateable_area[1] ),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.D(_0077_),
    .Q(\updateable_area[2] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.D(_0078_),
    .Q(\updateable_area[3] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.D(_0079_),
    .Q(\updateable_area[4] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.D(_0080_),
    .Q(\updateable_area[5] ),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.D(_0081_),
    .Q(\updateable_area[6] ),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.D(_0082_),
    .Q(\updateable_area[7] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.D(_0083_),
    .Q(\updateable_area[8] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.D(_0084_),
    .Q(\updateable_area[9] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.D(_0085_),
    .Q(\updateable_area[10] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.D(_0086_),
    .Q(\updateable_area[11] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.D(_0087_),
    .Q(\updateable_area[12] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.D(_0088_),
    .Q(\updateable_area[13] ),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.D(_0089_),
    .Q(\updateable_area[14] ),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.D(_0090_),
    .Q(\updateable_area[15] ),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.D(_0091_),
    .Q(\updateable_area[16] ),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.D(_0092_),
    .Q(\updateable_area[17] ),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.D(_0093_),
    .Q(\updateable_area[18] ),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.D(_0094_),
    .Q(\updateable_area[19] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.D(_0095_),
    .Q(\updateable_area[20] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.D(_0096_),
    .Q(\updateable_area[21] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.D(_0097_),
    .Q(\updateable_area[22] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.D(_0098_),
    .Q(\updateable_area[23] ),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.D(_0099_),
    .Q(\updateable_area[24] ),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.D(_0100_),
    .Q(\updateable_area[25] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.D(_0101_),
    .Q(\updateable_area[26] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.D(_0102_),
    .Q(\updateable_area[27] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.D(_0103_),
    .Q(\updateable_area[28] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.D(_0104_),
    .Q(\updateable_area[29] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.D(_0105_),
    .Q(\updateable_area[30] ),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.D(_0106_),
    .Q(\updateable_area[31] ),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.D(_0107_),
    .Q(\disruptive_area[0] ),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.D(_0108_),
    .Q(\disruptive_area[1] ),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.D(_0109_),
    .Q(\disruptive_area[2] ),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.D(_0110_),
    .Q(\disruptive_area[3] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.D(_0111_),
    .Q(\disruptive_area[4] ),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.D(_0112_),
    .Q(\disruptive_area[5] ),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.D(_0113_),
    .Q(\disruptive_area[6] ),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.D(_0114_),
    .Q(\disruptive_area[7] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.D(_0115_),
    .Q(\disruptive_area[8] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.D(_0116_),
    .Q(\disruptive_area[9] ),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.D(_0117_),
    .Q(\disruptive_area[10] ),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.D(_0118_),
    .Q(\disruptive_area[11] ),
    .CLK(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.D(_0119_),
    .Q(\disruptive_area[12] ),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.D(_0120_),
    .Q(\disruptive_area[13] ),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.D(_0121_),
    .Q(\disruptive_area[14] ),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.D(_0122_),
    .Q(\disruptive_area[15] ),
    .CLK(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.D(_0123_),
    .Q(\disruptive_area[16] ),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.D(_0124_),
    .Q(\disruptive_area[17] ),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.D(_0125_),
    .Q(\disruptive_area[18] ),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.D(_0126_),
    .Q(\disruptive_area[19] ),
    .CLK(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.D(_0127_),
    .Q(\disruptive_area[20] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.D(_0128_),
    .Q(\disruptive_area[21] ),
    .CLK(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.D(_0129_),
    .Q(\disruptive_area[22] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.D(_0130_),
    .Q(\disruptive_area[23] ),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.D(_0131_),
    .Q(\disruptive_area[24] ),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.D(_0132_),
    .Q(\disruptive_area[25] ),
    .CLK(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.D(_0133_),
    .Q(\disruptive_area[26] ),
    .CLK(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.D(_0134_),
    .Q(\disruptive_area[27] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.D(_0135_),
    .Q(\disruptive_area[28] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.D(_0136_),
    .Q(\disruptive_area[29] ),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.D(_0137_),
    .Q(\disruptive_area[30] ),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.D(_0138_),
    .Q(\disruptive_area[31] ),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.D(_0139_),
    .Q(net129),
    .CLK(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.D(_0140_),
    .Q(net140),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.D(_0141_),
    .Q(net151),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_2 _1190_ (.D(_0142_),
    .Q(net154),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.D(_0143_),
    .Q(net155),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.D(_0144_),
    .Q(net156),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.D(_0145_),
    .Q(net157),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.D(_0146_),
    .Q(net158),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.D(_0147_),
    .Q(net159),
    .CLK(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.D(_0148_),
    .Q(net160),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.D(_0149_),
    .Q(net130),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.D(_0150_),
    .Q(net131),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.D(_0151_),
    .Q(net132),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.D(_0152_),
    .Q(net133),
    .CLK(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.D(_0153_),
    .Q(net134),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.D(_0154_),
    .Q(net135),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.D(_0155_),
    .Q(net136),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.D(_0156_),
    .Q(net137),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.D(_0157_),
    .Q(net138),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.D(_0158_),
    .Q(net139),
    .CLK(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.D(_0159_),
    .Q(net141),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.D(_0160_),
    .Q(net142),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.D(_0161_),
    .Q(net143),
    .CLK(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.D(_0162_),
    .Q(net144),
    .CLK(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.D(_0163_),
    .Q(net145),
    .CLK(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.D(_0164_),
    .Q(net146),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.D(_0165_),
    .Q(net147),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.D(_0166_),
    .Q(net148),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.D(_0167_),
    .Q(net149),
    .CLK(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.D(_0168_),
    .Q(net150),
    .CLK(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.D(_0169_),
    .Q(net152),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.D(_0170_),
    .Q(net153),
    .CLK(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(i_copro_crm[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(i_copro_crm[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(i_copro_crm[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(i_copro_crm[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(i_copro_crn[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(i_copro_crn[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(i_copro_crn[2]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(i_copro_crn[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(i_copro_num[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(i_copro_num[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(i_copro_num[2]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(i_copro_num[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(i_copro_opcode1[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(i_copro_opcode1[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(i_copro_opcode1[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(i_copro_opcode2[0]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(i_copro_opcode2[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(i_copro_opcode2[2]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(i_copro_operation[0]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(i_copro_operation[1]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(i_copro_write_data[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(i_copro_write_data[10]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(i_copro_write_data[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(i_copro_write_data[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(i_copro_write_data[13]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(i_copro_write_data[14]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(i_copro_write_data[15]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(i_copro_write_data[16]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(i_copro_write_data[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(i_copro_write_data[18]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(i_copro_write_data[19]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(i_copro_write_data[1]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(i_copro_write_data[20]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(i_copro_write_data[21]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(i_copro_write_data[22]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(i_copro_write_data[23]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(i_copro_write_data[24]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(i_copro_write_data[25]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(i_copro_write_data[26]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(i_copro_write_data[27]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(i_copro_write_data[28]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(i_copro_write_data[29]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(i_copro_write_data[2]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(i_copro_write_data[30]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(i_copro_write_data[31]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(i_copro_write_data[3]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(i_copro_write_data[4]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(i_copro_write_data[5]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(i_copro_write_data[6]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(i_copro_write_data[7]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(i_copro_write_data[8]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(i_copro_write_data[9]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(i_core_stall),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(i_fault),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(i_fault_address[0]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(i_fault_address[10]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(i_fault_address[11]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(i_fault_address[12]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(i_fault_address[13]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(i_fault_address[14]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(i_fault_address[15]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(i_fault_address[16]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(i_fault_address[17]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(i_fault_address[18]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(i_fault_address[19]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(i_fault_address[1]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(i_fault_address[20]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(i_fault_address[21]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(i_fault_address[22]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(i_fault_address[23]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(i_fault_address[24]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(i_fault_address[25]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(i_fault_address[26]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(i_fault_address[27]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(i_fault_address[28]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(i_fault_address[29]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(i_fault_address[2]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(i_fault_address[30]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(i_fault_address[31]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(i_fault_address[3]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(i_fault_address[4]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(i_fault_address[5]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(i_fault_address[6]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(i_fault_address[7]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(i_fault_address[8]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(i_fault_address[9]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(i_fault_status[0]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(i_fault_status[1]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(i_fault_status[2]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(i_fault_status[3]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(i_fault_status[4]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(i_fault_status[5]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(i_fault_status[6]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(i_fault_status[7]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 output95 (.A(net95),
    .X(o_cache_enable));
 sky130_fd_sc_hd__clkbuf_2 output96 (.A(net96),
    .X(o_cache_flush));
 sky130_fd_sc_hd__clkbuf_2 output97 (.A(net97),
    .X(o_cacheable_area[0]));
 sky130_fd_sc_hd__clkbuf_2 output98 (.A(net98),
    .X(o_cacheable_area[10]));
 sky130_fd_sc_hd__clkbuf_2 output99 (.A(net99),
    .X(o_cacheable_area[11]));
 sky130_fd_sc_hd__clkbuf_2 output100 (.A(net100),
    .X(o_cacheable_area[12]));
 sky130_fd_sc_hd__clkbuf_2 output101 (.A(net101),
    .X(o_cacheable_area[13]));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(o_cacheable_area[14]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(o_cacheable_area[15]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(o_cacheable_area[16]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(o_cacheable_area[17]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(o_cacheable_area[18]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(o_cacheable_area[19]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(o_cacheable_area[1]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(o_cacheable_area[20]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(o_cacheable_area[21]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(o_cacheable_area[22]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(o_cacheable_area[23]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(o_cacheable_area[24]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(o_cacheable_area[25]));
 sky130_fd_sc_hd__clkbuf_2 output115 (.A(net115),
    .X(o_cacheable_area[26]));
 sky130_fd_sc_hd__clkbuf_2 output116 (.A(net116),
    .X(o_cacheable_area[27]));
 sky130_fd_sc_hd__clkbuf_2 output117 (.A(net117),
    .X(o_cacheable_area[28]));
 sky130_fd_sc_hd__clkbuf_2 output118 (.A(net118),
    .X(o_cacheable_area[29]));
 sky130_fd_sc_hd__clkbuf_2 output119 (.A(net119),
    .X(o_cacheable_area[2]));
 sky130_fd_sc_hd__clkbuf_2 output120 (.A(net120),
    .X(o_cacheable_area[30]));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(o_cacheable_area[31]));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(o_cacheable_area[3]));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(o_cacheable_area[4]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(o_cacheable_area[5]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(o_cacheable_area[6]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(o_cacheable_area[7]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(o_cacheable_area[8]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(o_cacheable_area[9]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(o_copro_read_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(o_copro_read_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(o_copro_read_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(o_copro_read_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(o_copro_read_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(o_copro_read_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(o_copro_read_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(o_copro_read_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(o_copro_read_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(o_copro_read_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(o_copro_read_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(o_copro_read_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(o_copro_read_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(o_copro_read_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(o_copro_read_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(o_copro_read_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(o_copro_read_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(o_copro_read_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(o_copro_read_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(o_copro_read_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(o_copro_read_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(o_copro_read_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(o_copro_read_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(o_copro_read_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(o_copro_read_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(o_copro_read_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(o_copro_read_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(o_copro_read_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(o_copro_read_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(o_copro_read_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(o_copro_read_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(o_copro_read_data[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_15_0_i_clk));
endmodule
