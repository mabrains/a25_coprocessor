* NGSPICE file created from a25_coprocessor.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt a25_coprocessor i_clk i_copro_crm[0] i_copro_crm[1] i_copro_crm[2] i_copro_crm[3]
+ i_copro_crn[0] i_copro_crn[1] i_copro_crn[2] i_copro_crn[3] i_copro_num[0] i_copro_num[1]
+ i_copro_num[2] i_copro_num[3] i_copro_opcode1[0] i_copro_opcode1[1] i_copro_opcode1[2]
+ i_copro_opcode2[0] i_copro_opcode2[1] i_copro_opcode2[2] i_copro_operation[0] i_copro_operation[1]
+ i_copro_write_data[0] i_copro_write_data[10] i_copro_write_data[11] i_copro_write_data[12]
+ i_copro_write_data[13] i_copro_write_data[14] i_copro_write_data[15] i_copro_write_data[16]
+ i_copro_write_data[17] i_copro_write_data[18] i_copro_write_data[19] i_copro_write_data[1]
+ i_copro_write_data[20] i_copro_write_data[21] i_copro_write_data[22] i_copro_write_data[23]
+ i_copro_write_data[24] i_copro_write_data[25] i_copro_write_data[26] i_copro_write_data[27]
+ i_copro_write_data[28] i_copro_write_data[29] i_copro_write_data[2] i_copro_write_data[30]
+ i_copro_write_data[31] i_copro_write_data[3] i_copro_write_data[4] i_copro_write_data[5]
+ i_copro_write_data[6] i_copro_write_data[7] i_copro_write_data[8] i_copro_write_data[9]
+ i_core_stall i_fault i_fault_address[0] i_fault_address[10] i_fault_address[11]
+ i_fault_address[12] i_fault_address[13] i_fault_address[14] i_fault_address[15]
+ i_fault_address[16] i_fault_address[17] i_fault_address[18] i_fault_address[19]
+ i_fault_address[1] i_fault_address[20] i_fault_address[21] i_fault_address[22] i_fault_address[23]
+ i_fault_address[24] i_fault_address[25] i_fault_address[26] i_fault_address[27]
+ i_fault_address[28] i_fault_address[29] i_fault_address[2] i_fault_address[30] i_fault_address[31]
+ i_fault_address[3] i_fault_address[4] i_fault_address[5] i_fault_address[6] i_fault_address[7]
+ i_fault_address[8] i_fault_address[9] i_fault_status[0] i_fault_status[1] i_fault_status[2]
+ i_fault_status[3] i_fault_status[4] i_fault_status[5] i_fault_status[6] i_fault_status[7]
+ o_cache_enable o_cache_flush o_cacheable_area[0] o_cacheable_area[10] o_cacheable_area[11]
+ o_cacheable_area[12] o_cacheable_area[13] o_cacheable_area[14] o_cacheable_area[15]
+ o_cacheable_area[16] o_cacheable_area[17] o_cacheable_area[18] o_cacheable_area[19]
+ o_cacheable_area[1] o_cacheable_area[20] o_cacheable_area[21] o_cacheable_area[22]
+ o_cacheable_area[23] o_cacheable_area[24] o_cacheable_area[25] o_cacheable_area[26]
+ o_cacheable_area[27] o_cacheable_area[28] o_cacheable_area[29] o_cacheable_area[2]
+ o_cacheable_area[30] o_cacheable_area[31] o_cacheable_area[3] o_cacheable_area[4]
+ o_cacheable_area[5] o_cacheable_area[6] o_cacheable_area[7] o_cacheable_area[8]
+ o_cacheable_area[9] o_copro_read_data[0] o_copro_read_data[10] o_copro_read_data[11]
+ o_copro_read_data[12] o_copro_read_data[13] o_copro_read_data[14] o_copro_read_data[15]
+ o_copro_read_data[16] o_copro_read_data[17] o_copro_read_data[18] o_copro_read_data[19]
+ o_copro_read_data[1] o_copro_read_data[20] o_copro_read_data[21] o_copro_read_data[22]
+ o_copro_read_data[23] o_copro_read_data[24] o_copro_read_data[25] o_copro_read_data[26]
+ o_copro_read_data[27] o_copro_read_data[28] o_copro_read_data[29] o_copro_read_data[2]
+ o_copro_read_data[30] o_copro_read_data[31] o_copro_read_data[3] o_copro_read_data[4]
+ o_copro_read_data[5] o_copro_read_data[6] o_copro_read_data[7] o_copro_read_data[8]
+ o_copro_read_data[9] VPWR VGND
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0985_ _0985_/A VGND VGND VPWR VPWR _0985_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0770_ _0993_/A _0993_/B _0944_/D VGND VGND VPWR VPWR _0770_/X sky130_fd_sc_hd__or3_4
X_1184_ _1215_/CLK _1184_/D VGND VGND VPWR VPWR _1184_/Q sky130_fd_sc_hd__dfxtp_1
X_0968_ _1077_/Q _0963_/X input30/X _0964_/X VGND VGND VPWR VPWR _1077_/D sky130_fd_sc_hd__a22o_1
X_0899_ _0927_/A VGND VGND VPWR VPWR _0899_/X sky130_fd_sc_hd__buf_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0822_ _1172_/Q _0816_/X input29/X _0817_/X VGND VGND VPWR VPWR _1172_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0684_ _1135_/Q VGND VGND VPWR VPWR _0684_/Y sky130_fd_sc_hd__inv_2
X_0753_ _1095_/Q VGND VGND VPWR VPWR _0753_/Y sky130_fd_sc_hd__inv_2
X_1098_ _1176_/CLK _1098_/D VGND VGND VPWR VPWR _1098_/Q sky130_fd_sc_hd__dfxtp_1
X_1167_ _1206_/CLK _1167_/D VGND VGND VPWR VPWR _1167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ _1065_/Q VGND VGND VPWR VPWR _1021_/X sky130_fd_sc_hd__buf_2
X_0805_ _1185_/Q _0800_/X input44/X _0803_/X VGND VGND VPWR VPWR _1185_/D sky130_fd_sc_hd__a22o_1
X_0667_ _1105_/Q VGND VGND VPWR VPWR _0667_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0736_ _0736_/A _1054_/Q VGND VGND VPWR VPWR _0736_/X sky130_fd_sc_hd__or2b_1
X_0598_ _0581_/X _1210_/Q _0572_/X _0597_/Y VGND VGND VPWR VPWR _1210_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ _0993_/A input6/X _0944_/D VGND VGND VPWR VPWR _0522_/A sky130_fd_sc_hd__or3_4
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1004_ _1050_/Q _1000_/X input89/X _1001_/X VGND VGND VPWR VPWR _1050_/D sky130_fd_sc_hd__a22o_1
X_0719_ _0704_/X _1195_/Q _0695_/X _0718_/Y VGND VGND VPWR VPWR _1195_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput97 _1059_/Q VGND VGND VPWR VPWR o_cacheable_area[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0984_ _0984_/A VGND VGND VPWR VPWR _0984_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1183_ _1215_/CLK _1183_/D VGND VGND VPWR VPWR _1183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0967_ _1078_/Q _0963_/X input31/X _0964_/X VGND VGND VPWR VPWR _1078_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0898_ _1001_/A VGND VGND VPWR VPWR _0927_/A sky130_fd_sc_hd__buf_2
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0821_ _1173_/Q _0816_/X input30/X _0817_/X VGND VGND VPWR VPWR _1173_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0752_ _1063_/Q VGND VGND VPWR VPWR _0752_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0683_ _1103_/Q VGND VGND VPWR VPWR _0683_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1166_ _1166_/CLK _1166_/D VGND VGND VPWR VPWR _1166_/Q sky130_fd_sc_hd__dfxtp_1
X_1097_ _1209_/CLK _1097_/D VGND VGND VPWR VPWR _1097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1020_ _1064_/Q VGND VGND VPWR VPWR _1020_/X sky130_fd_sc_hd__buf_2
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0735_ _1097_/Q VGND VGND VPWR VPWR _0735_/Y sky130_fd_sc_hd__inv_2
X_0804_ _1186_/Q _0800_/X input45/X _0803_/X VGND VGND VPWR VPWR _1186_/D sky130_fd_sc_hd__a22o_1
X_0666_ _0666_/A VGND VGND VPWR VPWR _0666_/X sky130_fd_sc_hd__clkbuf_4
X_0597_ _0590_/Y _0574_/X _0591_/Y _0592_/X _0596_/X VGND VGND VPWR VPWR _0597_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1149_ _1181_/CLK _1149_/D VGND VGND VPWR VPWR _1149_/Q sky130_fd_sc_hd__dfxtp_1
X_1218_ _1218_/CLK _1218_/D VGND VGND VPWR VPWR _1218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0520_ input8/X input7/X VGND VGND VPWR VPWR _0944_/D sky130_fd_sc_hd__or2_2
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1003_ _1051_/Q _1000_/X input90/X _1001_/X VGND VGND VPWR VPWR _1051_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0718_ _0713_/Y _0706_/X _0522_/A _0717_/X VGND VGND VPWR VPWR _0718_/Y sky130_fd_sc_hd__o211ai_2
X_0649_ _1107_/Q VGND VGND VPWR VPWR _0649_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput98 _1069_/Q VGND VGND VPWR VPWR o_cacheable_area[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_i_clk clkbuf_3_7_0_i_clk/X VGND VGND VPWR VPWR _1200_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0983_ _1066_/Q _0977_/X input50/X _0978_/X VGND VGND VPWR VPWR _1066_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1182_ _1215_/CLK _1182_/D VGND VGND VPWR VPWR _1182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0966_ _1079_/Q _0963_/X input33/X _0964_/X VGND VGND VPWR VPWR _1079_/D sky130_fd_sc_hd__a22o_1
X_0897_ _1000_/A VGND VGND VPWR VPWR _1001_/A sky130_fd_sc_hd__inv_2
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0820_ _1174_/Q _0816_/X input31/X _0817_/X VGND VGND VPWR VPWR _1174_/D sky130_fd_sc_hd__a22o_1
X_0751_ _1127_/Q VGND VGND VPWR VPWR _0751_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0682_ _1071_/Q VGND VGND VPWR VPWR _0682_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1165_ _1195_/CLK _1165_/D VGND VGND VPWR VPWR _1165_/Q sky130_fd_sc_hd__dfxtp_1
X_1096_ _1216_/CLK _1096_/D VGND VGND VPWR VPWR _1096_/Q sky130_fd_sc_hd__dfxtp_1
X_0949_ _0985_/A VGND VGND VPWR VPWR _0964_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0665_ _1073_/Q VGND VGND VPWR VPWR _0665_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0734_ _1065_/Q VGND VGND VPWR VPWR _0734_/Y sky130_fd_sc_hd__inv_2
X_0803_ _0817_/A VGND VGND VPWR VPWR _0803_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0596_ _0593_/Y _0594_/X _0595_/Y _0554_/X VGND VGND VPWR VPWR _0596_/X sky130_fd_sc_hd__o22a_1
X_1079_ _1174_/CLK _1079_/D VGND VGND VPWR VPWR _1079_/Q sky130_fd_sc_hd__dfxtp_2
X_1148_ _1181_/CLK _1148_/D VGND VGND VPWR VPWR _1148_/Q sky130_fd_sc_hd__dfxtp_1
X_1217_ _1218_/CLK _1217_/D VGND VGND VPWR VPWR _1217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_i_clk clkbuf_3_5_0_i_clk/X VGND VGND VPWR VPWR _1210_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1002_ _1052_/Q _1000_/X input91/X _1001_/X VGND VGND VPWR VPWR _1052_/D sky130_fd_sc_hd__a22o_1
X_0717_ _0714_/Y _0617_/X _0715_/Y _0619_/X _0716_/X VGND VGND VPWR VPWR _0717_/X
+ sky130_fd_sc_hd__o221a_1
X_0648_ _1075_/Q VGND VGND VPWR VPWR _0648_/Y sky130_fd_sc_hd__inv_2
X_0579_ _0573_/Y _0574_/X _0575_/Y _0541_/X _0578_/X VGND VGND VPWR VPWR _0579_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput99 _1070_/Q VGND VGND VPWR VPWR o_cacheable_area[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0982_ _1067_/Q _0977_/X input51/X _0978_/X VGND VGND VPWR VPWR _1067_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1181_ _1181_/CLK _1181_/D VGND VGND VPWR VPWR _1181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0965_ _1080_/Q _0963_/X input34/X _0964_/X VGND VGND VPWR VPWR _1080_/D sky130_fd_sc_hd__a22o_1
X_0896_ _0926_/A VGND VGND VPWR VPWR _0896_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0681_ _1167_/Q VGND VGND VPWR VPWR _0681_/Y sky130_fd_sc_hd__inv_2
X_0750_ _1159_/Q VGND VGND VPWR VPWR _0750_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1164_ _1211_/CLK _1164_/D VGND VGND VPWR VPWR _1164_/Q sky130_fd_sc_hd__dfxtp_1
X_1095_ _1216_/CLK _1095_/D VGND VGND VPWR VPWR _1095_/Q sky130_fd_sc_hd__dfxtp_1
X_0948_ _0984_/A VGND VGND VPWR VPWR _0985_/A sky130_fd_sc_hd__inv_2
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0879_ _0886_/A VGND VGND VPWR VPWR _0879_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0802_ _0838_/A VGND VGND VPWR VPWR _0817_/A sky130_fd_sc_hd__clkbuf_2
X_0664_ _1169_/Q VGND VGND VPWR VPWR _0664_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0733_ _1129_/Q VGND VGND VPWR VPWR _0733_/Y sky130_fd_sc_hd__inv_2
X_1216_ _1216_/CLK _1216_/D VGND VGND VPWR VPWR _1216_/Q sky130_fd_sc_hd__dfxtp_1
X_0595_ _1146_/Q VGND VGND VPWR VPWR _0595_/Y sky130_fd_sc_hd__inv_2
X_1078_ _1211_/CLK _1078_/D VGND VGND VPWR VPWR _1078_/Q sky130_fd_sc_hd__dfxtp_2
X_1147_ _1180_/CLK _1147_/D VGND VGND VPWR VPWR _1147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1001_ _1001_/A VGND VGND VPWR VPWR _1001_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0716_ _0716_/A _1099_/Q VGND VGND VPWR VPWR _0716_/X sky130_fd_sc_hd__or2b_1
X_0647_ _1171_/Q VGND VGND VPWR VPWR _0647_/Y sky130_fd_sc_hd__inv_2
X_0578_ _0576_/Y _0544_/X _0577_/Y _0554_/X VGND VGND VPWR VPWR _0578_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_i_clk clkbuf_4_9_0_i_clk/A VGND VGND VPWR VPWR _1187_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0981_ _1068_/Q _0977_/X input52/X _0978_/X VGND VGND VPWR VPWR _1068_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1180_ _1180_/CLK _1180_/D VGND VGND VPWR VPWR _1180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0964_ _0964_/A VGND VGND VPWR VPWR _0964_/X sky130_fd_sc_hd__clkbuf_2
X_0895_ _1000_/A VGND VGND VPWR VPWR _0926_/A sky130_fd_sc_hd__buf_2
Xclkbuf_3_6_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_3_6_0_i_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0680_ _0663_/X _1200_/Q _0654_/X _0679_/Y VGND VGND VPWR VPWR _1200_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1163_ _1166_/CLK _1163_/D VGND VGND VPWR VPWR _1163_/Q sky130_fd_sc_hd__dfxtp_1
X_1094_ _1209_/CLK _1094_/D VGND VGND VPWR VPWR _1094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0947_ _0963_/A VGND VGND VPWR VPWR _0947_/X sky130_fd_sc_hd__clkbuf_2
X_0878_ _0885_/A VGND VGND VPWR VPWR _0878_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0801_ _0837_/A VGND VGND VPWR VPWR _0838_/A sky130_fd_sc_hd__inv_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0594_ _0668_/A VGND VGND VPWR VPWR _0594_/X sky130_fd_sc_hd__clkbuf_2
X_0663_ _0798_/A VGND VGND VPWR VPWR _0663_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0732_ _1161_/Q VGND VGND VPWR VPWR _0732_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1215_ _1215_/CLK _1215_/D VGND VGND VPWR VPWR _1215_/Q sky130_fd_sc_hd__dfxtp_1
X_1146_ _1180_/CLK _1146_/D VGND VGND VPWR VPWR _1146_/Q sky130_fd_sc_hd__dfxtp_1
X_1077_ _1174_/CLK _1077_/D VGND VGND VPWR VPWR _1077_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1000_ _1000_/A VGND VGND VPWR VPWR _1000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0715_ _1163_/Q VGND VGND VPWR VPWR _0715_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_5_0_i_clk clkbuf_4_5_0_i_clk/A VGND VGND VPWR VPWR _1176_/CLK sky130_fd_sc_hd__clkbuf_1
X_0646_ _0625_/X _1204_/Q _0614_/X _0645_/Y VGND VGND VPWR VPWR _1204_/D sky130_fd_sc_hd__a22o_1
X_0577_ _1148_/Q VGND VGND VPWR VPWR _0577_/Y sky130_fd_sc_hd__inv_2
X_1129_ _1187_/CLK _1129_/D VGND VGND VPWR VPWR _1129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0629_ _1142_/Q VGND VGND VPWR VPWR _0629_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_i_clk i_clk VGND VGND VPWR VPWR clkbuf_0_i_clk/X sky130_fd_sc_hd__clkbuf_16
X_0980_ _1069_/Q _0977_/X input22/X _0978_/X VGND VGND VPWR VPWR _1069_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_4_5_0_i_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0963_ _0963_/A VGND VGND VPWR VPWR _0963_/X sky130_fd_sc_hd__clkbuf_2
X_0894_ _0894_/A _0894_/B VGND VGND VPWR VPWR _1000_/A sky130_fd_sc_hd__nand2_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1162_ _1195_/CLK _1162_/D VGND VGND VPWR VPWR _1162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1093_ _1216_/CLK _1093_/D VGND VGND VPWR VPWR _1093_/Q sky130_fd_sc_hd__dfxtp_1
X_0877_ _1135_/Q _0871_/X input24/X _0872_/X VGND VGND VPWR VPWR _1135_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0946_ _0984_/A VGND VGND VPWR VPWR _0963_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0731_ _0704_/X _1194_/Q _0695_/X _0730_/Y VGND VGND VPWR VPWR _1194_/D sky130_fd_sc_hd__a22o_1
X_0800_ _0816_/A VGND VGND VPWR VPWR _0800_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0662_ _0625_/X _1202_/Q _0654_/X _0661_/Y VGND VGND VPWR VPWR _1202_/D sky130_fd_sc_hd__a22o_1
X_0593_ _1114_/Q VGND VGND VPWR VPWR _0593_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1214_ _1215_/CLK _1214_/D VGND VGND VPWR VPWR _1214_/Q sky130_fd_sc_hd__dfxtp_1
X_1145_ _1181_/CLK _1145_/D VGND VGND VPWR VPWR _1145_/Q sky130_fd_sc_hd__dfxtp_1
X_1076_ _1174_/CLK _1076_/D VGND VGND VPWR VPWR _1076_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_1_0_i_clk clkbuf_4_1_0_i_clk/A VGND VGND VPWR VPWR _1180_/CLK sky130_fd_sc_hd__clkbuf_1
X_0929_ _1101_/Q _0926_/X input56/X _0927_/X VGND VGND VPWR VPWR _1101_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0714_ _1067_/Q VGND VGND VPWR VPWR _0714_/Y sky130_fd_sc_hd__inv_2
X_0645_ _0640_/Y _0583_/X _0522_/A _0644_/X VGND VGND VPWR VPWR _0645_/Y sky130_fd_sc_hd__o211ai_1
X_0576_ _1116_/Q VGND VGND VPWR VPWR _0576_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1128_ _1210_/CLK _1128_/D VGND VGND VPWR VPWR _1128_/Q sky130_fd_sc_hd__dfxtp_1
X_1059_ _1187_/CLK _1059_/D VGND VGND VPWR VPWR _1059_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0628_ _1110_/Q VGND VGND VPWR VPWR _0628_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0559_ _1086_/Q VGND VGND VPWR VPWR _0559_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0962_ _1081_/Q _0956_/X input35/X _0957_/X VGND VGND VPWR VPWR _1081_/D sky130_fd_sc_hd__a22o_1
X_0893_ _1123_/Q _0864_/A input21/X _0865_/A VGND VGND VPWR VPWR _1123_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1092_ _1216_/CLK _1092_/D VGND VGND VPWR VPWR _1092_/Q sky130_fd_sc_hd__dfxtp_1
X_1161_ _1187_/CLK _1161_/D VGND VGND VPWR VPWR _1161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0876_ _1136_/Q _0871_/X input25/X _0872_/X VGND VGND VPWR VPWR _1136_/D sky130_fd_sc_hd__a22o_1
X_0945_ _1007_/A _0993_/B _1007_/C VGND VGND VPWR VPWR _0984_/A sky130_fd_sc_hd__or3_4
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0730_ _0720_/Y _0697_/X _0721_/Y _0706_/X _0729_/X VGND VGND VPWR VPWR _0730_/Y
+ sky130_fd_sc_hd__o221ai_2
X_0661_ _0655_/Y _0656_/X _0657_/Y _0592_/X _0660_/X VGND VGND VPWR VPWR _0661_/Y
+ sky130_fd_sc_hd__o221ai_2
X_0592_ _0666_/A VGND VGND VPWR VPWR _0592_/X sky130_fd_sc_hd__buf_4
X_1213_ _1215_/CLK _1213_/D VGND VGND VPWR VPWR _1213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ _1176_/CLK _1144_/D VGND VGND VPWR VPWR _1144_/Q sky130_fd_sc_hd__dfxtp_1
X_1075_ _1206_/CLK _1075_/D VGND VGND VPWR VPWR _1075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ _1102_/Q _0926_/X input57/X _0927_/X VGND VGND VPWR VPWR _1102_/D sky130_fd_sc_hd__a22o_1
X_0859_ _1149_/Q _0857_/X input39/X _0858_/X VGND VGND VPWR VPWR _1149_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0713_ _1131_/Q VGND VGND VPWR VPWR _0713_/Y sky130_fd_sc_hd__inv_2
X_0644_ _0641_/Y _0617_/X _0642_/Y _0619_/X _0643_/X VGND VGND VPWR VPWR _0644_/X
+ sky130_fd_sc_hd__o221a_1
X_0575_ _1084_/Q VGND VGND VPWR VPWR _0575_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1058_ _1187_/CLK _1058_/D VGND VGND VPWR VPWR _1058_/Q sky130_fd_sc_hd__dfxtp_1
X_1127_ _1209_/CLK _1127_/D VGND VGND VPWR VPWR _1127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0627_ _1078_/Q VGND VGND VPWR VPWR _0627_/Y sky130_fd_sc_hd__inv_2
X_0558_ _1182_/Q VGND VGND VPWR VPWR _0558_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0961_ _1082_/Q _0956_/X input36/X _0957_/X VGND VGND VPWR VPWR _1082_/D sky130_fd_sc_hd__a22o_1
X_0892_ _1124_/Q _0864_/A input32/X _0865_/A VGND VGND VPWR VPWR _1124_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1091_ _1216_/CLK _1091_/D VGND VGND VPWR VPWR _1091_/Q sky130_fd_sc_hd__dfxtp_1
X_1160_ _1210_/CLK _1160_/D VGND VGND VPWR VPWR _1160_/Q sky130_fd_sc_hd__dfxtp_1
X_0944_ _0944_/A _0944_/B _0944_/C _0944_/D VGND VGND VPWR VPWR _1007_/C sky130_fd_sc_hd__or4_4
X_0875_ _1137_/Q _0871_/X input26/X _0872_/X VGND VGND VPWR VPWR _1137_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0660_ _0658_/Y _0594_/X _0659_/Y _0610_/X VGND VGND VPWR VPWR _0660_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0591_ _1082_/Q VGND VGND VPWR VPWR _0591_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1212_ _1215_/CLK _1212_/D VGND VGND VPWR VPWR _1212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1074_ _1170_/CLK _1074_/D VGND VGND VPWR VPWR _1074_/Q sky130_fd_sc_hd__dfxtp_2
X_1143_ _1176_/CLK _1143_/D VGND VGND VPWR VPWR _1143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0927_ _0927_/A VGND VGND VPWR VPWR _0927_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0789_ _1091_/Q VGND VGND VPWR VPWR _0789_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0858_ _0865_/A VGND VGND VPWR VPWR _0858_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0643_ _0716_/A _1108_/Q VGND VGND VPWR VPWR _0643_/X sky130_fd_sc_hd__or2b_1
X_0574_ _0697_/A VGND VGND VPWR VPWR _0574_/X sky130_fd_sc_hd__buf_4
X_0712_ _0704_/X _1196_/Q _0695_/X _0711_/Y VGND VGND VPWR VPWR _1196_/D sky130_fd_sc_hd__a22o_1
X_1126_ _1209_/CLK _1126_/D VGND VGND VPWR VPWR _1126_/Q sky130_fd_sc_hd__dfxtp_1
X_1057_ _1170_/CLK _1057_/D VGND VGND VPWR VPWR _1057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0626_ _1174_/Q VGND VGND VPWR VPWR _0626_/Y sky130_fd_sc_hd__inv_2
X_0557_ _0537_/X _1215_/Q _0511_/X _0556_/Y VGND VGND VPWR VPWR _1215_/D sky130_fd_sc_hd__a22o_1
X_1109_ _1176_/CLK _1109_/D VGND VGND VPWR VPWR _1109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0609_ _1144_/Q VGND VGND VPWR VPWR _0609_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0960_ _1083_/Q _0956_/X input37/X _0957_/X VGND VGND VPWR VPWR _1083_/D sky130_fd_sc_hd__a22o_1
X_0891_ _1125_/Q _0885_/X input43/X _0886_/X VGND VGND VPWR VPWR _1125_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1090_ _1218_/CLK _1090_/D VGND VGND VPWR VPWR _1090_/Q sky130_fd_sc_hd__dfxtp_2
X_0874_ _1138_/Q _0871_/X input27/X _0872_/X VGND VGND VPWR VPWR _1138_/D sky130_fd_sc_hd__a22o_1
X_0943_ _1091_/Q _0940_/X input55/X _0941_/X VGND VGND VPWR VPWR _1091_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0590_ _1178_/Q VGND VGND VPWR VPWR _0590_/Y sky130_fd_sc_hd__inv_2
X_1142_ _1176_/CLK _1142_/D VGND VGND VPWR VPWR _1142_/Q sky130_fd_sc_hd__dfxtp_1
X_1211_ _1211_/CLK _1211_/D VGND VGND VPWR VPWR _1211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1073_ _1200_/CLK _1073_/D VGND VGND VPWR VPWR _1073_/Q sky130_fd_sc_hd__dfxtp_2
X_0926_ _0926_/A VGND VGND VPWR VPWR _0926_/X sky130_fd_sc_hd__clkbuf_2
X_0857_ _0864_/A VGND VGND VPWR VPWR _0857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0788_ _1123_/Q VGND VGND VPWR VPWR _0788_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0711_ _0705_/Y _0706_/X _0522_/A _0710_/X VGND VGND VPWR VPWR _0711_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0642_ _1172_/Q VGND VGND VPWR VPWR _0642_/Y sky130_fd_sc_hd__inv_2
X_0573_ _1180_/Q VGND VGND VPWR VPWR _0573_/Y sky130_fd_sc_hd__inv_2
X_1125_ _1209_/CLK _1125_/D VGND VGND VPWR VPWR _1125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ _1170_/CLK _1056_/D VGND VGND VPWR VPWR _1056_/Q sky130_fd_sc_hd__dfxtp_2
X_0909_ _1115_/Q _0905_/X input71/X _0906_/X VGND VGND VPWR VPWR _1115_/D sky130_fd_sc_hd__a22o_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0625_ _0625_/A VGND VGND VPWR VPWR _0625_/X sky130_fd_sc_hd__clkbuf_2
X_0556_ _0550_/Y _0518_/X _0551_/Y _0541_/X _0555_/X VGND VGND VPWR VPWR _0556_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1108_ _1176_/CLK _1108_/D VGND VGND VPWR VPWR _1108_/Q sky130_fd_sc_hd__dfxtp_1
X_1039_ _1083_/Q VGND VGND VPWR VPWR _1039_/X sky130_fd_sc_hd__buf_2
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0608_ _1112_/Q VGND VGND VPWR VPWR _0608_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0539_ _1088_/Q VGND VGND VPWR VPWR _0539_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0890_ _1126_/Q _0885_/X input46/X _0886_/X VGND VGND VPWR VPWR _1126_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0873_ _1139_/Q _0871_/X input28/X _0872_/X VGND VGND VPWR VPWR _1139_/D sky130_fd_sc_hd__a22o_1
X_0942_ _1092_/Q _0940_/X input66/X _0941_/X VGND VGND VPWR VPWR _1092_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1072_ _1200_/CLK _1072_/D VGND VGND VPWR VPWR _1072_/Q sky130_fd_sc_hd__dfxtp_1
X_1210_ _1210_/CLK _1210_/D VGND VGND VPWR VPWR _1210_/Q sky130_fd_sc_hd__dfxtp_1
X_1141_ _1174_/CLK _1141_/D VGND VGND VPWR VPWR _1141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0925_ _1103_/Q _0919_/X input58/X _0920_/X VGND VGND VPWR VPWR _1103_/D sky130_fd_sc_hd__a22o_1
X_0856_ _1150_/Q _0848_/X input40/X _0851_/X VGND VGND VPWR VPWR _1150_/D sky130_fd_sc_hd__a22o_1
X_0787_ _1059_/Q VGND VGND VPWR VPWR _0787_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0710_ _0707_/Y _0617_/X _0708_/Y _0619_/X _0709_/X VGND VGND VPWR VPWR _0710_/X
+ sky130_fd_sc_hd__o221a_1
X_0641_ _1076_/Q VGND VGND VPWR VPWR _0641_/Y sky130_fd_sc_hd__inv_2
X_0572_ _0614_/A VGND VGND VPWR VPWR _0572_/X sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1055_ _1216_/CLK _1055_/D VGND VGND VPWR VPWR _1055_/Q sky130_fd_sc_hd__dfxtp_1
X_1124_ _1211_/CLK _1124_/D VGND VGND VPWR VPWR _1124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0908_ _1116_/Q _0905_/X input72/X _0906_/X VGND VGND VPWR VPWR _1116_/D sky130_fd_sc_hd__a22o_1
X_0839_ _1161_/Q _0837_/X input49/X _0838_/X VGND VGND VPWR VPWR _1161_/D sky130_fd_sc_hd__a22o_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0624_ _0581_/X _1207_/Q _0614_/X _0623_/Y VGND VGND VPWR VPWR _1207_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0555_ _0552_/Y _0544_/X _0553_/Y _0554_/X VGND VGND VPWR VPWR _0555_/X sky130_fd_sc_hd__o22a_1
X_1107_ _1195_/CLK _1107_/D VGND VGND VPWR VPWR _1107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1038_ _1082_/Q VGND VGND VPWR VPWR _1038_/X sky130_fd_sc_hd__buf_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0607_ _1080_/Q VGND VGND VPWR VPWR _0607_/Y sky130_fd_sc_hd__inv_2
X_0538_ _1184_/Q VGND VGND VPWR VPWR _0538_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0941_ _1001_/A VGND VGND VPWR VPWR _0941_/X sky130_fd_sc_hd__clkbuf_2
X_0872_ _0886_/A VGND VGND VPWR VPWR _0872_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ _1195_/CLK _1071_/D VGND VGND VPWR VPWR _1071_/Q sky130_fd_sc_hd__dfxtp_2
X_1140_ _1174_/CLK _1140_/D VGND VGND VPWR VPWR _1140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0924_ _1104_/Q _0919_/X input59/X _0920_/X VGND VGND VPWR VPWR _1104_/D sky130_fd_sc_hd__a22o_1
X_0855_ _1151_/Q _0848_/X input41/X _0851_/X VGND VGND VPWR VPWR _1151_/D sky130_fd_sc_hd__a22o_1
X_0786_ _0749_/X _1188_/Q _0740_/X _0785_/Y VGND VGND VPWR VPWR _1188_/D sky130_fd_sc_hd__a22o_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0640_ _1140_/Q VGND VGND VPWR VPWR _0640_/Y sky130_fd_sc_hd__inv_2
X_0571_ _0537_/X _1213_/Q _0511_/X _0570_/Y VGND VGND VPWR VPWR _1213_/D sky130_fd_sc_hd__a22o_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1054_ _1216_/CLK _1054_/D VGND VGND VPWR VPWR _1054_/Q sky130_fd_sc_hd__dfxtp_1
X_1123_ _1187_/CLK _1123_/D VGND VGND VPWR VPWR _1123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0907_ _1117_/Q _0905_/X input73/X _0906_/X VGND VGND VPWR VPWR _1117_/D sky130_fd_sc_hd__a22o_1
X_0769_ _1058_/Q VGND VGND VPWR VPWR _0769_/Y sky130_fd_sc_hd__inv_2
X_0838_ _0838_/A VGND VGND VPWR VPWR _0838_/X sky130_fd_sc_hd__clkbuf_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0623_ _0615_/Y _0583_/X _0522_/X _0622_/X VGND VGND VPWR VPWR _0623_/Y sky130_fd_sc_hd__o211ai_4
X_0554_ _0706_/A VGND VGND VPWR VPWR _0554_/X sky130_fd_sc_hd__clkbuf_2
X_1106_ _1195_/CLK _1106_/D VGND VGND VPWR VPWR _1106_/Q sky130_fd_sc_hd__dfxtp_1
X_1037_ _1081_/Q VGND VGND VPWR VPWR _1037_/X sky130_fd_sc_hd__buf_2
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput90 i_fault_status[3] VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_1
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_i_clk clkbuf_3_7_0_i_clk/X VGND VGND VPWR VPWR _1206_/CLK sky130_fd_sc_hd__clkbuf_1
X_0606_ _1176_/Q VGND VGND VPWR VPWR _0606_/Y sky130_fd_sc_hd__inv_2
X_0537_ _0625_/A VGND VGND VPWR VPWR _0537_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0940_ _1000_/A VGND VGND VPWR VPWR _0940_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0871_ _0885_/A VGND VGND VPWR VPWR _0871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1070_ _1166_/CLK _1070_/D VGND VGND VPWR VPWR _1070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0923_ _1105_/Q _0919_/X input60/X _0920_/X VGND VGND VPWR VPWR _1105_/D sky130_fd_sc_hd__a22o_1
X_0854_ _1152_/Q _0848_/X input42/X _0851_/X VGND VGND VPWR VPWR _1152_/D sky130_fd_sc_hd__a22o_1
X_0785_ _0777_/Y _0736_/A _0778_/Y _0541_/A _0784_/X VGND VGND VPWR VPWR _0785_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1199_ _1200_/CLK _1199_/D VGND VGND VPWR VPWR _1199_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0570_ _0565_/Y _0518_/X _0566_/Y _0541_/X _0569_/X VGND VGND VPWR VPWR _0570_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1122_ _1211_/CLK _1122_/D VGND VGND VPWR VPWR _1122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1053_ _1216_/CLK _1053_/D VGND VGND VPWR VPWR _1053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0906_ _0927_/A VGND VGND VPWR VPWR _0906_/X sky130_fd_sc_hd__clkbuf_2
X_0837_ _0837_/A VGND VGND VPWR VPWR _0837_/X sky130_fd_sc_hd__clkbuf_2
X_0699_ _1101_/Q VGND VGND VPWR VPWR _0699_/Y sky130_fd_sc_hd__inv_2
X_0768_ _1125_/Q VGND VGND VPWR VPWR _0768_/Y sky130_fd_sc_hd__inv_2
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_i_clk clkbuf_3_5_0_i_clk/X VGND VGND VPWR VPWR _1209_/CLK sky130_fd_sc_hd__clkbuf_1
X_0622_ _0616_/Y _0617_/X _0618_/Y _0619_/X _0621_/X VGND VGND VPWR VPWR _0622_/X
+ sky130_fd_sc_hd__o221a_1
X_0553_ _1151_/Q VGND VGND VPWR VPWR _0553_/Y sky130_fd_sc_hd__inv_2
X_1105_ _1200_/CLK _1105_/D VGND VGND VPWR VPWR _1105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1036_ _1080_/Q VGND VGND VPWR VPWR _1036_/X sky130_fd_sc_hd__buf_2
Xinput80 i_fault_address[3] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_1
Xinput91 i_fault_status[4] VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0536_ _1217_/Q _0625_/A _0511_/X _0535_/Y VGND VGND VPWR VPWR _1217_/D sky130_fd_sc_hd__a22o_1
X_0605_ _0581_/X _1209_/Q _0572_/X _0604_/Y VGND VGND VPWR VPWR _1209_/D sky130_fd_sc_hd__a22o_1
X_1019_ _1063_/Q VGND VGND VPWR VPWR _1019_/X sky130_fd_sc_hd__buf_2
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0519_ input5/X VGND VGND VPWR VPWR _0993_/A sky130_fd_sc_hd__buf_1
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0870_ _1140_/Q _0864_/X input29/X _0865_/X VGND VGND VPWR VPWR _1140_/D sky130_fd_sc_hd__a22o_1
X_0999_ _1053_/Q _0940_/X input92/X _0941_/X VGND VGND VPWR VPWR _1053_/D sky130_fd_sc_hd__a22o_1
XFILLER_10_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0922_ _1106_/Q _0919_/X input61/X _0920_/X VGND VGND VPWR VPWR _1106_/D sky130_fd_sc_hd__a22o_1
X_0853_ _1153_/Q _0848_/X input44/X _0851_/X VGND VGND VPWR VPWR _1153_/D sky130_fd_sc_hd__a22o_1
X_0784_ _0779_/Y _0706_/A _0780_/Y _0770_/X _0783_/X VGND VGND VPWR VPWR _0784_/X
+ sky130_fd_sc_hd__o221a_1
Xinput1 i_copro_crm[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_1
X_1198_ _1200_/CLK _1198_/D VGND VGND VPWR VPWR _1198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1052_ _1209_/CLK _1052_/D VGND VGND VPWR VPWR _1052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ _1180_/CLK _1121_/D VGND VGND VPWR VPWR _1121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0836_ _1162_/Q _0830_/X input50/X _0831_/X VGND VGND VPWR VPWR _1162_/D sky130_fd_sc_hd__a22o_1
X_0905_ _0926_/A VGND VGND VPWR VPWR _0905_/X sky130_fd_sc_hd__clkbuf_2
X_0767_ _1061_/Q VGND VGND VPWR VPWR _0767_/Y sky130_fd_sc_hd__inv_2
X_0698_ _1069_/Q VGND VGND VPWR VPWR _0698_/Y sky130_fd_sc_hd__inv_2
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0621_ _0716_/A _1111_/Q VGND VGND VPWR VPWR _0621_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0552_ _1119_/Q VGND VGND VPWR VPWR _0552_/Y sky130_fd_sc_hd__inv_2
X_1104_ _1195_/CLK _1104_/D VGND VGND VPWR VPWR _1104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1035_ _1079_/Q VGND VGND VPWR VPWR _1035_/X sky130_fd_sc_hd__buf_2
X_0819_ _1175_/Q _0816_/X input33/X _0817_/X VGND VGND VPWR VPWR _1175_/D sky130_fd_sc_hd__a22o_1
Xinput92 i_fault_status[5] VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_1
Xinput81 i_fault_address[4] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_1
Xinput70 i_fault_address[23] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0604_ _0599_/Y _0583_/X _0522_/X _0603_/X VGND VGND VPWR VPWR _0604_/Y sky130_fd_sc_hd__o211ai_4
Xclkbuf_4_8_0_i_clk clkbuf_4_9_0_i_clk/A VGND VGND VPWR VPWR _1216_/CLK sky130_fd_sc_hd__clkbuf_1
X_0535_ _0512_/Y _0518_/X _0522_/X _0534_/X VGND VGND VPWR VPWR _0535_/Y sky130_fd_sc_hd__o211ai_1
X_1018_ _1062_/Q VGND VGND VPWR VPWR _1018_/X sky130_fd_sc_hd__buf_2
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0518_ _0518_/A VGND VGND VPWR VPWR _0518_/X sky130_fd_sc_hd__buf_2
XFILLER_49_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0998_ _1054_/Q _0940_/X input93/X _0941_/X VGND VGND VPWR VPWR _1054_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_3_5_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_3_5_0_i_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0921_ _1107_/Q _0919_/X input62/X _0920_/X VGND VGND VPWR VPWR _1107_/D sky130_fd_sc_hd__a22o_1
X_0852_ _1154_/Q _0848_/X input45/X _0851_/X VGND VGND VPWR VPWR _1154_/D sky130_fd_sc_hd__a22o_1
X_0783_ _0781_/Y _0668_/A _0782_/Y _0798_/D VGND VGND VPWR VPWR _0783_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1197_ _1200_/CLK _1197_/D VGND VGND VPWR VPWR _1197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 i_copro_crm[1] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_1
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ _1209_/CLK _1051_/D VGND VGND VPWR VPWR _1051_/Q sky130_fd_sc_hd__dfxtp_1
X_1120_ _1215_/CLK _1120_/D VGND VGND VPWR VPWR _1120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0904_ _1118_/Q _0896_/X input74/X _0899_/X VGND VGND VPWR VPWR _1118_/D sky130_fd_sc_hd__a22o_1
X_0835_ _1163_/Q _0830_/X input51/X _0831_/X VGND VGND VPWR VPWR _1163_/D sky130_fd_sc_hd__a22o_1
X_0697_ _0697_/A VGND VGND VPWR VPWR _0697_/X sky130_fd_sc_hd__clkbuf_4
X_0766_ _1050_/Q VGND VGND VPWR VPWR _0766_/Y sky130_fd_sc_hd__inv_2
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0620_ _0725_/A VGND VGND VPWR VPWR _0716_/A sky130_fd_sc_hd__buf_1
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0551_ _1087_/Q VGND VGND VPWR VPWR _0551_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1034_ _1078_/Q VGND VGND VPWR VPWR _1034_/X sky130_fd_sc_hd__buf_2
X_1103_ _1200_/CLK _1103_/D VGND VGND VPWR VPWR _1103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_4_0_i_clk clkbuf_4_5_0_i_clk/A VGND VGND VPWR VPWR _1174_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0818_ _1176_/Q _0816_/X input34/X _0817_/X VGND VGND VPWR VPWR _1176_/D sky130_fd_sc_hd__a22o_1
Xinput93 i_fault_status[6] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_1
Xinput82 i_fault_address[5] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_1
Xinput71 i_fault_address[24] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_1
Xinput60 i_fault_address[14] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_1
X_0749_ _0798_/A VGND VGND VPWR VPWR _0749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0603_ _0600_/Y _0666_/A _0601_/Y _0518_/A _0602_/X VGND VGND VPWR VPWR _0603_/X
+ sky130_fd_sc_hd__o221a_1
X_0534_ _0523_/Y _0666_/A _0528_/Y _0706_/A _0533_/X VGND VGND VPWR VPWR _0534_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1017_ _1061_/Q VGND VGND VPWR VPWR _1017_/X sky130_fd_sc_hd__buf_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0517_ _0697_/A VGND VGND VPWR VPWR _0518_/A sky130_fd_sc_hd__buf_2
Xclkbuf_3_1_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_4_3_0_i_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0997_ _1055_/Q _0940_/X input94/X _0941_/X VGND VGND VPWR VPWR _1055_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0920_ _0927_/A VGND VGND VPWR VPWR _0920_/X sky130_fd_sc_hd__clkbuf_2
X_0851_ _0865_/A VGND VGND VPWR VPWR _0851_/X sky130_fd_sc_hd__clkbuf_2
X_0782_ _1156_/Q VGND VGND VPWR VPWR _0782_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1196_ _1206_/CLK _1196_/D VGND VGND VPWR VPWR _1196_/Q sky130_fd_sc_hd__dfxtp_1
Xinput3 i_copro_crm[2] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_1
XFILLER_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1050_ _1209_/CLK _1050_/D VGND VGND VPWR VPWR _1050_/Q sky130_fd_sc_hd__dfxtp_1
X_0834_ _1164_/Q _0830_/X input52/X _0831_/X VGND VGND VPWR VPWR _1164_/D sky130_fd_sc_hd__a22o_1
X_0903_ _1119_/Q _0896_/X input75/X _0899_/X VGND VGND VPWR VPWR _1119_/D sky130_fd_sc_hd__a22o_1
X_0696_ _1165_/Q VGND VGND VPWR VPWR _0696_/Y sky130_fd_sc_hd__inv_2
X_0765_ _0749_/X _1190_/Q _0740_/X _0764_/Y VGND VGND VPWR VPWR _1190_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_4_0_0_i_clk clkbuf_4_1_0_i_clk/A VGND VGND VPWR VPWR _1181_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1179_ _1180_/CLK _1179_/D VGND VGND VPWR VPWR _1179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0550_ _1183_/Q VGND VGND VPWR VPWR _0550_/Y sky130_fd_sc_hd__inv_2
X_1102_ _1176_/CLK _1102_/D VGND VGND VPWR VPWR _1102_/Q sky130_fd_sc_hd__dfxtp_1
X_1033_ _1077_/Q VGND VGND VPWR VPWR _1033_/X sky130_fd_sc_hd__buf_2
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput50 i_copro_write_data[7] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_2
Xinput61 i_fault_address[15] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_1
Xinput72 i_fault_address[25] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_1
X_0817_ _0817_/A VGND VGND VPWR VPWR _0817_/X sky130_fd_sc_hd__clkbuf_2
X_0679_ _0673_/Y _0656_/X _0674_/Y _0666_/X _0678_/X VGND VGND VPWR VPWR _0679_/Y
+ sky130_fd_sc_hd__o221ai_1
Xinput83 i_fault_address[6] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_1
Xinput94 i_fault_status[7] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__buf_1
X_0748_ _0704_/X _1192_/Q _0740_/X _0747_/Y VGND VGND VPWR VPWR _1192_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0602_ _0602_/A _1113_/Q VGND VGND VPWR VPWR _0602_/X sky130_fd_sc_hd__or2b_1
X_0533_ _0602_/A _1121_/Q VGND VGND VPWR VPWR _0533_/X sky130_fd_sc_hd__or2b_1
X_1016_ _1060_/Q VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__buf_2
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0516_ _0798_/D VGND VGND VPWR VPWR _0697_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0996_ input21/X _1056_/Q _0996_/S VGND VGND VPWR VPWR _1056_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0850_ _0886_/A VGND VGND VPWR VPWR _0865_/A sky130_fd_sc_hd__clkbuf_2
X_0781_ _1092_/Q VGND VGND VPWR VPWR _0781_/Y sky130_fd_sc_hd__inv_2
Xinput4 i_copro_crm[3] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1195_ _1195_/CLK _1195_/D VGND VGND VPWR VPWR _1195_/Q sky130_fd_sc_hd__dfxtp_1
X_0979_ _1070_/Q _0977_/X input23/X _0978_/X VGND VGND VPWR VPWR _1070_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0833_ _1165_/Q _0830_/X input22/X _0831_/X VGND VGND VPWR VPWR _1165_/D sky130_fd_sc_hd__a22o_1
X_0902_ _1120_/Q _0896_/X input76/X _0899_/X VGND VGND VPWR VPWR _1120_/D sky130_fd_sc_hd__a22o_1
X_0764_ _0758_/Y _0518_/A _0759_/Y _0583_/A _0763_/X VGND VGND VPWR VPWR _0764_/Y
+ sky130_fd_sc_hd__o221ai_2
X_0695_ _0894_/A VGND VGND VPWR VPWR _0695_/X sky130_fd_sc_hd__clkbuf_2
X_1178_ _1180_/CLK _1178_/D VGND VGND VPWR VPWR _1178_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput160 _1196_/Q VGND VGND VPWR VPWR o_copro_read_data[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1101_ _1176_/CLK _1101_/D VGND VGND VPWR VPWR _1101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1032_ _1076_/Q VGND VGND VPWR VPWR _1032_/X sky130_fd_sc_hd__buf_2
XFILLER_23_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput62 i_fault_address[16] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
Xinput84 i_fault_address[7] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_1
Xinput40 i_copro_write_data[27] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_2
X_0816_ _0816_/A VGND VGND VPWR VPWR _0816_/X sky130_fd_sc_hd__clkbuf_2
Xinput73 i_fault_address[26] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__buf_1
Xinput51 i_copro_write_data[8] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
X_0747_ _0741_/Y _0697_/X _0742_/Y _0706_/X _0746_/X VGND VGND VPWR VPWR _0747_/Y
+ sky130_fd_sc_hd__o221ai_2
X_0678_ _0675_/Y _0668_/X _0676_/Y _0677_/X VGND VGND VPWR VPWR _0678_/X sky130_fd_sc_hd__o22a_1
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0601_ _1177_/Q VGND VGND VPWR VPWR _0601_/Y sky130_fd_sc_hd__inv_2
X_0532_ _0725_/A VGND VGND VPWR VPWR _0602_/A sky130_fd_sc_hd__buf_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1015_ _1059_/Q VGND VGND VPWR VPWR _1015_/X sky130_fd_sc_hd__buf_2
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0515_ input8/X _0726_/B _1007_/A input6/X VGND VGND VPWR VPWR _0798_/D sky130_fd_sc_hd__or4_4
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0995_ input32/X _1057_/Q _0996_/S VGND VGND VPWR VPWR _1057_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0780_ _1057_/Q VGND VGND VPWR VPWR _0780_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 i_copro_crn[0] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_1
X_1194_ _1200_/CLK _1194_/D VGND VGND VPWR VPWR _1194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0978_ _0985_/A VGND VGND VPWR VPWR _0978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0832_ _1166_/Q _0830_/X input23/X _0831_/X VGND VGND VPWR VPWR _1166_/D sky130_fd_sc_hd__a22o_1
X_0763_ _0760_/Y _0723_/X _0761_/Y _0602_/A _0762_/X VGND VGND VPWR VPWR _0763_/X
+ sky130_fd_sc_hd__o221a_1
X_0901_ _1121_/Q _0896_/X input78/X _0899_/X VGND VGND VPWR VPWR _1121_/D sky130_fd_sc_hd__a22o_1
X_0694_ _0663_/X _1198_/Q _0654_/X _0693_/Y VGND VGND VPWR VPWR _1198_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1177_ _1181_/CLK _1177_/D VGND VGND VPWR VPWR _1177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 _1216_/Q VGND VGND VPWR VPWR o_copro_read_data[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1100_ _1176_/CLK _1100_/D VGND VGND VPWR VPWR _1100_/Q sky130_fd_sc_hd__dfxtp_1
X_1031_ _1075_/Q VGND VGND VPWR VPWR _1031_/X sky130_fd_sc_hd__buf_2
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput41 i_copro_write_data[28] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_2
Xinput74 i_fault_address[27] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__buf_1
Xinput85 i_fault_address[8] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_1
Xinput52 i_copro_write_data[9] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
Xinput30 i_copro_write_data[18] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_2
Xinput63 i_fault_address[17] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_2
X_0746_ _0743_/Y _0723_/X _0744_/Y _0725_/X _0745_/X VGND VGND VPWR VPWR _0746_/X
+ sky130_fd_sc_hd__o221a_1
X_0815_ _1177_/Q _0809_/X input35/X _0810_/X VGND VGND VPWR VPWR _1177_/D sky130_fd_sc_hd__a22o_1
X_0677_ _0846_/D VGND VGND VPWR VPWR _0677_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0531_ _1007_/A _0993_/B input8/X _0726_/B VGND VGND VPWR VPWR _0725_/A sky130_fd_sc_hd__or4_4
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0600_ _1081_/Q VGND VGND VPWR VPWR _0600_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1014_ _0625_/A _1218_/Q _0614_/A _1013_/Y VGND VGND VPWR VPWR _1218_/D sky130_fd_sc_hd__a22o_1
X_0729_ _0722_/Y _0723_/X _0724_/Y _0725_/X _0728_/X VGND VGND VPWR VPWR _0729_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_43_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0514_ input5/X VGND VGND VPWR VPWR _1007_/A sky130_fd_sc_hd__inv_2
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ input43/X _1058_/Q _0996_/S VGND VGND VPWR VPWR _1058_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 i_copro_crn[1] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_2
X_1193_ _1210_/CLK _1193_/D VGND VGND VPWR VPWR _1193_/Q sky130_fd_sc_hd__dfxtp_1
X_0977_ _0984_/A VGND VGND VPWR VPWR _0977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0900_ _1122_/Q _0896_/X input79/X _0899_/X VGND VGND VPWR VPWR _1122_/D sky130_fd_sc_hd__a22o_1
X_0693_ _0688_/Y _0656_/X _0689_/Y _0666_/X _0692_/X VGND VGND VPWR VPWR _0693_/Y
+ sky130_fd_sc_hd__o221ai_4
X_0831_ _0838_/A VGND VGND VPWR VPWR _0831_/X sky130_fd_sc_hd__clkbuf_2
X_0762_ _0762_/A _1051_/Q VGND VGND VPWR VPWR _0762_/X sky130_fd_sc_hd__or2b_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1176_ _1176_/CLK _1176_/D VGND VGND VPWR VPWR _1176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput151 _1189_/Q VGND VGND VPWR VPWR o_copro_read_data[2] sky130_fd_sc_hd__clkbuf_2
Xoutput140 _1188_/Q VGND VGND VPWR VPWR o_copro_read_data[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1030_ _1074_/Q VGND VGND VPWR VPWR _1030_/X sky130_fd_sc_hd__buf_2
Xinput20 i_copro_operation[1] VGND VGND VPWR VPWR _0797_/A sky130_fd_sc_hd__buf_1
Xinput31 i_copro_write_data[19] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0814_ _1178_/Q _0809_/X input36/X _0810_/X VGND VGND VPWR VPWR _1178_/D sky130_fd_sc_hd__a22o_1
Xinput64 i_fault_address[18] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
X_0676_ _1136_/Q VGND VGND VPWR VPWR _0676_/Y sky130_fd_sc_hd__inv_2
Xinput42 i_copro_write_data[29] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_2
Xinput75 i_fault_address[28] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_1
Xinput86 i_fault_address[9] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_1
Xinput53 i_core_stall VGND VGND VPWR VPWR _0944_/A sky130_fd_sc_hd__buf_2
X_0745_ _0762_/A _1053_/Q VGND VGND VPWR VPWR _0745_/X sky130_fd_sc_hd__or2b_1
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1159_ _1209_/CLK _1159_/D VGND VGND VPWR VPWR _1159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0530_ _0846_/D VGND VGND VPWR VPWR _0706_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1013_ _1008_/Y _0518_/A _1009_/Y _0541_/A _1012_/X VGND VGND VPWR VPWR _1013_/Y
+ sky130_fd_sc_hd__o221ai_2
X_0659_ _1138_/Q VGND VGND VPWR VPWR _0659_/Y sky130_fd_sc_hd__inv_2
X_0728_ _0736_/A _1055_/Q VGND VGND VPWR VPWR _0728_/X sky130_fd_sc_hd__or2b_1
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0513_ input7/X VGND VGND VPWR VPWR _0726_/B sky130_fd_sc_hd__inv_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0993_ _0993_/A _0993_/B _1007_/C VGND VGND VPWR VPWR _0996_/S sky130_fd_sc_hd__or3_4
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 i_copro_crn[2] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_2
X_1192_ _1206_/CLK _1192_/D VGND VGND VPWR VPWR _1192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0976_ _1071_/Q _0970_/X input24/X _0971_/X VGND VGND VPWR VPWR _1071_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ _0837_/A VGND VGND VPWR VPWR _0830_/X sky130_fd_sc_hd__clkbuf_2
X_0692_ _0690_/Y _0668_/X _0691_/Y _0677_/X VGND VGND VPWR VPWR _0692_/X sky130_fd_sc_hd__o22a_1
X_0761_ _1094_/Q VGND VGND VPWR VPWR _0761_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1175_ _1176_/CLK _1175_/D VGND VGND VPWR VPWR _1175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0959_ _1084_/Q _0956_/X input38/X _0957_/X VGND VGND VPWR VPWR _1084_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput141 _1207_/Q VGND VGND VPWR VPWR o_copro_read_data[20] sky130_fd_sc_hd__clkbuf_2
Xoutput152 _1217_/Q VGND VGND VPWR VPWR o_copro_read_data[30] sky130_fd_sc_hd__clkbuf_2
Xoutput130 _1197_/Q VGND VGND VPWR VPWR o_copro_read_data[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 i_copro_write_data[1] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_2
Xinput21 i_copro_write_data[0] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_2
Xinput43 i_copro_write_data[2] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput10 i_copro_num[1] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_1
X_0813_ _1179_/Q _0809_/X input37/X _0810_/X VGND VGND VPWR VPWR _1179_/D sky130_fd_sc_hd__a22o_1
Xinput54 i_fault VGND VGND VPWR VPWR _0894_/B sky130_fd_sc_hd__buf_1
X_0675_ _1104_/Q VGND VGND VPWR VPWR _0675_/Y sky130_fd_sc_hd__inv_2
Xinput76 i_fault_address[29] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__clkbuf_1
X_0744_ _1096_/Q VGND VGND VPWR VPWR _0744_/Y sky130_fd_sc_hd__inv_2
Xinput87 i_fault_status[0] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__clkbuf_1
Xinput65 i_fault_address[19] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1158_ _1209_/CLK _1158_/D VGND VGND VPWR VPWR _1158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1089_ _1218_/CLK _1089_/D VGND VGND VPWR VPWR _1089_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1012_ _1010_/Y _0725_/X _1011_/Y _0677_/X VGND VGND VPWR VPWR _1012_/X sky130_fd_sc_hd__o22a_1
X_0727_ _0762_/A VGND VGND VPWR VPWR _0736_/A sky130_fd_sc_hd__clkbuf_2
X_0658_ _1106_/Q VGND VGND VPWR VPWR _0658_/Y sky130_fd_sc_hd__inv_2
X_0589_ _0581_/X _1211_/Q _0572_/X _0588_/Y VGND VGND VPWR VPWR _1211_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0512_ _1185_/Q VGND VGND VPWR VPWR _0512_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0992_ _1059_/Q _0963_/A input21/X _0964_/A VGND VGND VPWR VPWR _1059_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 i_copro_crn[3] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
X_1191_ _1210_/CLK _1191_/D VGND VGND VPWR VPWR _1191_/Q sky130_fd_sc_hd__dfxtp_1
X_0975_ _1072_/Q _0970_/X input25/X _0971_/X VGND VGND VPWR VPWR _1072_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ _1062_/Q VGND VGND VPWR VPWR _0760_/Y sky130_fd_sc_hd__inv_2
X_0691_ _1134_/Q VGND VGND VPWR VPWR _0691_/Y sky130_fd_sc_hd__inv_2
X_1174_ _1174_/CLK _1174_/D VGND VGND VPWR VPWR _1174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0889_ _1127_/Q _0885_/X input47/X _0886_/X VGND VGND VPWR VPWR _1127_/D sky130_fd_sc_hd__a22o_1
X_0958_ _1085_/Q _0956_/X input39/X _0957_/X VGND VGND VPWR VPWR _1085_/D sky130_fd_sc_hd__a22o_1
Xoutput131 _1198_/Q VGND VGND VPWR VPWR o_copro_read_data[11] sky130_fd_sc_hd__clkbuf_2
Xoutput153 _1218_/Q VGND VGND VPWR VPWR o_copro_read_data[31] sky130_fd_sc_hd__clkbuf_2
Xoutput142 _1208_/Q VGND VGND VPWR VPWR o_copro_read_data[21] sky130_fd_sc_hd__clkbuf_2
Xoutput120 _1089_/Q VGND VGND VPWR VPWR o_cacheable_area[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput33 i_copro_write_data[20] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_2
Xinput22 i_copro_write_data[10] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_1
Xinput11 i_copro_num[2] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_1
Xinput66 i_fault_address[1] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_1
Xinput88 i_fault_status[1] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__clkbuf_1
Xinput77 i_fault_address[2] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
X_0743_ _1064_/Q VGND VGND VPWR VPWR _0743_/Y sky130_fd_sc_hd__inv_2
X_0812_ _1180_/Q _0809_/X input38/X _0810_/X VGND VGND VPWR VPWR _1180_/D sky130_fd_sc_hd__a22o_1
Xinput44 i_copro_write_data[30] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_1
Xinput55 i_fault_address[0] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_1
X_0674_ _1072_/Q VGND VGND VPWR VPWR _0674_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1157_ _1187_/CLK _1157_/D VGND VGND VPWR VPWR _1157_/Q sky130_fd_sc_hd__dfxtp_1
X_1088_ _1215_/CLK _1088_/D VGND VGND VPWR VPWR _1088_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1011_ _1154_/Q VGND VGND VPWR VPWR _1011_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0726_ input8/X _0726_/B _0993_/A _0726_/D VGND VGND VPWR VPWR _0762_/A sky130_fd_sc_hd__or4_4
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0657_ _1074_/Q VGND VGND VPWR VPWR _0657_/Y sky130_fd_sc_hd__inv_2
X_0588_ _0582_/Y _0583_/X _0522_/X _0587_/X VGND VGND VPWR VPWR _0588_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1209_ _1209_/CLK _1209_/D VGND VGND VPWR VPWR _1209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13_0_i_clk clkbuf_3_6_0_i_clk/X VGND VGND VPWR VPWR _1195_/CLK sky130_fd_sc_hd__clkbuf_1
X_0511_ _0614_/A VGND VGND VPWR VPWR _0511_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0709_ _0716_/A _1100_/Q VGND VGND VPWR VPWR _0709_/X sky130_fd_sc_hd__or2b_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0991_ _1060_/Q _0963_/A input32/X _0964_/A VGND VGND VPWR VPWR _1060_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 i_copro_num[0] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_1
XFILLER_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1190_ _1210_/CLK _1190_/D VGND VGND VPWR VPWR _1190_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0974_ _1073_/Q _0970_/X input26/X _0971_/X VGND VGND VPWR VPWR _1073_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0690_ _1102_/Q VGND VGND VPWR VPWR _0690_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1173_ _1174_/CLK _1173_/D VGND VGND VPWR VPWR _1173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput110 _1080_/Q VGND VGND VPWR VPWR o_cacheable_area[21] sky130_fd_sc_hd__clkbuf_2
Xoutput132 _1199_/Q VGND VGND VPWR VPWR o_copro_read_data[12] sky130_fd_sc_hd__clkbuf_2
Xoutput121 _1090_/Q VGND VGND VPWR VPWR o_cacheable_area[31] sky130_fd_sc_hd__clkbuf_2
Xoutput143 _1209_/Q VGND VGND VPWR VPWR o_copro_read_data[22] sky130_fd_sc_hd__clkbuf_2
X_0888_ _1128_/Q _0885_/X input48/X _0886_/X VGND VGND VPWR VPWR _1128_/D sky130_fd_sc_hd__a22o_1
X_0957_ _0964_/A VGND VGND VPWR VPWR _0957_/X sky130_fd_sc_hd__clkbuf_2
Xoutput154 _1190_/Q VGND VGND VPWR VPWR o_copro_read_data[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput34 i_copro_write_data[21] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_2
Xinput23 i_copro_write_data[11] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__buf_1
Xinput89 i_fault_status[2] VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_1
Xinput56 i_fault_address[10] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_1
Xinput67 i_fault_address[20] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__clkbuf_1
X_0673_ _1168_/Q VGND VGND VPWR VPWR _0673_/Y sky130_fd_sc_hd__inv_2
Xinput78 i_fault_address[30] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_1
Xinput12 i_copro_num[3] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_1
Xinput45 i_copro_write_data[31] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_2
X_0811_ _1181_/Q _0809_/X input39/X _0810_/X VGND VGND VPWR VPWR _1181_/D sky130_fd_sc_hd__a22o_1
X_0742_ _1128_/Q VGND VGND VPWR VPWR _0742_/Y sky130_fd_sc_hd__inv_2
X_1156_ _1170_/CLK _1156_/D VGND VGND VPWR VPWR _1156_/Q sky130_fd_sc_hd__dfxtp_1
X_1087_ _1218_/CLK _1087_/D VGND VGND VPWR VPWR _1087_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1010_ _1122_/Q VGND VGND VPWR VPWR _1010_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0725_ _0725_/A VGND VGND VPWR VPWR _0725_/X sky130_fd_sc_hd__buf_2
X_0656_ _0697_/A VGND VGND VPWR VPWR _0656_/X sky130_fd_sc_hd__clkbuf_4
X_1208_ _1210_/CLK _1208_/D VGND VGND VPWR VPWR _1208_/Q sky130_fd_sc_hd__dfxtp_1
X_0587_ _0584_/Y _0666_/A _0585_/Y _0518_/A _0586_/X VGND VGND VPWR VPWR _0587_/X
+ sky130_fd_sc_hd__o221a_1
X_1139_ _1170_/CLK _1139_/D VGND VGND VPWR VPWR _1139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0510_ _0894_/A VGND VGND VPWR VPWR _0614_/A sky130_fd_sc_hd__buf_1
X_0708_ _1164_/Q VGND VGND VPWR VPWR _0708_/Y sky130_fd_sc_hd__inv_2
X_0639_ _0625_/X _1205_/Q _0614_/X _0638_/Y VGND VGND VPWR VPWR _1205_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0990_ _1061_/Q _0984_/X input43/X _0985_/X VGND VGND VPWR VPWR _1061_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ _1074_/Q _0970_/X input27/X _0971_/X VGND VGND VPWR VPWR _1074_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1172_ _1174_/CLK _1172_/D VGND VGND VPWR VPWR _1172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ _0963_/A VGND VGND VPWR VPWR _0956_/X sky130_fd_sc_hd__clkbuf_2
Xoutput122 _1062_/Q VGND VGND VPWR VPWR o_cacheable_area[3] sky130_fd_sc_hd__clkbuf_2
Xoutput144 _1210_/Q VGND VGND VPWR VPWR o_copro_read_data[23] sky130_fd_sc_hd__clkbuf_2
Xoutput133 _1200_/Q VGND VGND VPWR VPWR o_copro_read_data[13] sky130_fd_sc_hd__clkbuf_2
Xoutput155 _1191_/Q VGND VGND VPWR VPWR o_copro_read_data[4] sky130_fd_sc_hd__clkbuf_2
Xoutput100 _1071_/Q VGND VGND VPWR VPWR o_cacheable_area[12] sky130_fd_sc_hd__clkbuf_2
Xoutput111 _1081_/Q VGND VGND VPWR VPWR o_cacheable_area[22] sky130_fd_sc_hd__clkbuf_2
X_0887_ _1129_/Q _0885_/X input49/X _0886_/X VGND VGND VPWR VPWR _1129_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 i_copro_opcode1[0] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_1
X_0810_ _0817_/A VGND VGND VPWR VPWR _0810_/X sky130_fd_sc_hd__clkbuf_2
Xinput79 i_fault_address[31] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__clkbuf_2
Xinput68 i_fault_address[21] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__buf_1
X_0672_ _0663_/X _1201_/Q _0654_/X _0671_/Y VGND VGND VPWR VPWR _1201_/D sky130_fd_sc_hd__a22o_1
Xinput46 i_copro_write_data[3] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_2
Xinput24 i_copro_write_data[12] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_2
Xinput57 i_fault_address[11] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_1
Xinput35 i_copro_write_data[22] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__buf_1
X_0741_ _1160_/Q VGND VGND VPWR VPWR _0741_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1086_ _1215_/CLK _1086_/D VGND VGND VPWR VPWR _1086_/Q sky130_fd_sc_hd__dfxtp_1
X_1155_ _1218_/CLK _1155_/D VGND VGND VPWR VPWR _1155_/Q sky130_fd_sc_hd__dfxtp_1
X_0939_ _1093_/Q _0933_/X input77/X _0934_/X VGND VGND VPWR VPWR _1093_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0724_ _1098_/Q VGND VGND VPWR VPWR _0724_/Y sky130_fd_sc_hd__inv_2
X_0655_ _1170_/Q VGND VGND VPWR VPWR _0655_/Y sky130_fd_sc_hd__inv_2
X_0586_ _0602_/A _1115_/Q VGND VGND VPWR VPWR _0586_/X sky130_fd_sc_hd__or2b_1
X_1207_ _1210_/CLK _1207_/D VGND VGND VPWR VPWR _1207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1069_ _1195_/CLK _1069_/D VGND VGND VPWR VPWR _1069_/Q sky130_fd_sc_hd__dfxtp_2
X_1138_ _1170_/CLK _1138_/D VGND VGND VPWR VPWR _1138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0707_ _1068_/Q VGND VGND VPWR VPWR _0707_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_7_0_i_clk clkbuf_4_7_0_i_clk/A VGND VGND VPWR VPWR _1166_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0569_ _0567_/Y _0544_/X _0568_/Y _0554_/X VGND VGND VPWR VPWR _0569_/X sky130_fd_sc_hd__o22a_1
X_0638_ _0633_/Y _0583_/X _0522_/X _0637_/X VGND VGND VPWR VPWR _0638_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ _1075_/Q _0970_/X input28/X _0971_/X VGND VGND VPWR VPWR _1075_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_4_9_0_i_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1171_ _1206_/CLK _1171_/D VGND VGND VPWR VPWR _1171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0955_ _1086_/Q _0947_/X input40/X _0950_/X VGND VGND VPWR VPWR _1086_/D sky130_fd_sc_hd__a22o_1
X_0886_ _0886_/A VGND VGND VPWR VPWR _0886_/X sky130_fd_sc_hd__clkbuf_2
Xoutput123 _1063_/Q VGND VGND VPWR VPWR o_cacheable_area[4] sky130_fd_sc_hd__clkbuf_2
Xoutput145 _1211_/Q VGND VGND VPWR VPWR o_copro_read_data[24] sky130_fd_sc_hd__clkbuf_2
Xoutput156 _1192_/Q VGND VGND VPWR VPWR o_copro_read_data[5] sky130_fd_sc_hd__clkbuf_2
Xoutput134 _1201_/Q VGND VGND VPWR VPWR o_copro_read_data[14] sky130_fd_sc_hd__clkbuf_2
Xoutput101 _1072_/Q VGND VGND VPWR VPWR o_cacheable_area[13] sky130_fd_sc_hd__clkbuf_2
Xoutput112 _1082_/Q VGND VGND VPWR VPWR o_cacheable_area[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput36 i_copro_write_data[23] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_2
Xinput25 i_copro_write_data[13] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_2
Xinput14 i_copro_opcode1[1] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_1
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0740_ _0894_/A VGND VGND VPWR VPWR _0740_/X sky130_fd_sc_hd__clkbuf_2
X_0671_ _0664_/Y _0656_/X _0665_/Y _0666_/X _0670_/X VGND VGND VPWR VPWR _0671_/Y
+ sky130_fd_sc_hd__o221ai_2
Xinput58 i_fault_address[12] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_1
Xinput69 i_fault_address[22] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
Xinput47 i_copro_write_data[4] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1154_ _1218_/CLK _1154_/D VGND VGND VPWR VPWR _1154_/Q sky130_fd_sc_hd__dfxtp_1
X_1085_ _1174_/CLK _1085_/D VGND VGND VPWR VPWR _1085_/Q sky130_fd_sc_hd__dfxtp_2
X_0938_ _1094_/Q _0933_/X input80/X _0934_/X VGND VGND VPWR VPWR _1094_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0869_ _1141_/Q _0864_/X input30/X _0865_/X VGND VGND VPWR VPWR _1141_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0723_ _0723_/A VGND VGND VPWR VPWR _0723_/X sky130_fd_sc_hd__buf_2
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0585_ _1179_/Q VGND VGND VPWR VPWR _0585_/Y sky130_fd_sc_hd__inv_2
X_0654_ _0894_/A VGND VGND VPWR VPWR _0654_/X sky130_fd_sc_hd__clkbuf_2
X_1137_ _1200_/CLK _1137_/D VGND VGND VPWR VPWR _1137_/Q sky130_fd_sc_hd__dfxtp_1
X_1206_ _1206_/CLK _1206_/D VGND VGND VPWR VPWR _1206_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_3_0_i_clk clkbuf_4_3_0_i_clk/A VGND VGND VPWR VPWR _1218_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1068_ _1166_/CLK _1068_/D VGND VGND VPWR VPWR _1068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0706_ _0706_/A VGND VGND VPWR VPWR _0706_/X sky130_fd_sc_hd__clkbuf_4
X_0637_ _0634_/Y _0617_/X _0635_/Y _0619_/X _0636_/X VGND VGND VPWR VPWR _0637_/X
+ sky130_fd_sc_hd__o221a_1
X_0568_ _1149_/Q VGND VGND VPWR VPWR _0568_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_4_1_0_i_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ _0985_/A VGND VGND VPWR VPWR _0971_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _1170_/CLK _1170_/D VGND VGND VPWR VPWR _1170_/Q sky130_fd_sc_hd__dfxtp_1
X_0954_ _1087_/Q _0947_/X input41/X _0950_/X VGND VGND VPWR VPWR _1087_/D sky130_fd_sc_hd__a22o_1
X_0885_ _0885_/A VGND VGND VPWR VPWR _0885_/X sky130_fd_sc_hd__clkbuf_2
Xoutput102 _1073_/Q VGND VGND VPWR VPWR o_cacheable_area[14] sky130_fd_sc_hd__clkbuf_2
Xoutput124 _1064_/Q VGND VGND VPWR VPWR o_cacheable_area[5] sky130_fd_sc_hd__clkbuf_2
Xoutput113 _1083_/Q VGND VGND VPWR VPWR o_cacheable_area[24] sky130_fd_sc_hd__clkbuf_2
Xoutput146 _1212_/Q VGND VGND VPWR VPWR o_copro_read_data[25] sky130_fd_sc_hd__clkbuf_2
Xoutput135 _1202_/Q VGND VGND VPWR VPWR o_copro_read_data[15] sky130_fd_sc_hd__clkbuf_2
Xoutput157 _1193_/Q VGND VGND VPWR VPWR o_copro_read_data[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 i_copro_write_data[14] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__buf_1
Xinput59 i_fault_address[13] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_1
X_0670_ _0667_/Y _0668_/X _0669_/Y _0610_/X VGND VGND VPWR VPWR _0670_/X sky130_fd_sc_hd__o22a_1
Xinput37 i_copro_write_data[24] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_1
Xinput48 i_copro_write_data[5] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_1
Xinput15 i_copro_opcode1[2] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_1
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1084_ _1181_/CLK _1084_/D VGND VGND VPWR VPWR _1084_/Q sky130_fd_sc_hd__dfxtp_1
X_1153_ _1218_/CLK _1153_/D VGND VGND VPWR VPWR _1153_/Q sky130_fd_sc_hd__dfxtp_1
X_0868_ _1142_/Q _0864_/X input31/X _0865_/X VGND VGND VPWR VPWR _1142_/D sky130_fd_sc_hd__a22o_1
X_0799_ _0837_/A VGND VGND VPWR VPWR _0816_/A sky130_fd_sc_hd__clkbuf_2
X_0937_ _1095_/Q _0933_/X input81/X _0934_/X VGND VGND VPWR VPWR _1095_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0722_ _1066_/Q VGND VGND VPWR VPWR _0722_/Y sky130_fd_sc_hd__inv_2
X_0653_ _0625_/X _1203_/Q _0614_/X _0652_/Y VGND VGND VPWR VPWR _1203_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0584_ _1083_/Q VGND VGND VPWR VPWR _0584_/Y sky130_fd_sc_hd__inv_2
X_1067_ _1166_/CLK _1067_/D VGND VGND VPWR VPWR _1067_/Q sky130_fd_sc_hd__dfxtp_1
X_1136_ _1200_/CLK _1136_/D VGND VGND VPWR VPWR _1136_/Q sky130_fd_sc_hd__dfxtp_1
X_1205_ _1206_/CLK _1205_/D VGND VGND VPWR VPWR _1205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0636_ _0716_/A _1109_/Q VGND VGND VPWR VPWR _0636_/X sky130_fd_sc_hd__or2b_1
X_0705_ _1132_/Q VGND VGND VPWR VPWR _0705_/Y sky130_fd_sc_hd__inv_2
X_0567_ _1117_/Q VGND VGND VPWR VPWR _0567_/Y sky130_fd_sc_hd__inv_2
X_1119_ _1215_/CLK _1119_/D VGND VGND VPWR VPWR _1119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0619_ _0798_/D VGND VGND VPWR VPWR _0619_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0970_ _0984_/A VGND VGND VPWR VPWR _0970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput125 _1065_/Q VGND VGND VPWR VPWR o_cacheable_area[6] sky130_fd_sc_hd__clkbuf_2
Xoutput103 _1074_/Q VGND VGND VPWR VPWR o_cacheable_area[15] sky130_fd_sc_hd__clkbuf_2
X_0884_ _1130_/Q _0878_/X input50/X _0879_/X VGND VGND VPWR VPWR _1130_/D sky130_fd_sc_hd__a22o_1
Xoutput114 _1084_/Q VGND VGND VPWR VPWR o_cacheable_area[25] sky130_fd_sc_hd__clkbuf_2
X_0953_ _1088_/Q _0947_/X input42/X _0950_/X VGND VGND VPWR VPWR _1088_/D sky130_fd_sc_hd__a22o_1
Xoutput158 _1194_/Q VGND VGND VPWR VPWR o_copro_read_data[7] sky130_fd_sc_hd__clkbuf_2
Xoutput136 _1203_/Q VGND VGND VPWR VPWR o_copro_read_data[16] sky130_fd_sc_hd__clkbuf_2
Xoutput147 _1213_/Q VGND VGND VPWR VPWR o_copro_read_data[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput16 i_copro_opcode2[0] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_1
Xinput38 i_copro_write_data[25] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_1
Xinput49 i_copro_write_data[6] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
Xinput27 i_copro_write_data[15] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__buf_2
X_1152_ _1215_/CLK _1152_/D VGND VGND VPWR VPWR _1152_/Q sky130_fd_sc_hd__dfxtp_1
X_1083_ _1180_/CLK _1083_/D VGND VGND VPWR VPWR _1083_/Q sky130_fd_sc_hd__dfxtp_1
X_0936_ _1096_/Q _0933_/X input82/X _0934_/X VGND VGND VPWR VPWR _1096_/D sky130_fd_sc_hd__a22o_1
X_0798_ _0798_/A _0944_/B _0944_/C _0798_/D VGND VGND VPWR VPWR _0837_/A sky130_fd_sc_hd__or4_4
X_0867_ _1143_/Q _0864_/X input33/X _0865_/X VGND VGND VPWR VPWR _1143_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0721_ _1130_/Q VGND VGND VPWR VPWR _0721_/Y sky130_fd_sc_hd__inv_2
X_0652_ _0647_/Y _0574_/X _0648_/Y _0592_/X _0651_/X VGND VGND VPWR VPWR _0652_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0583_ _0583_/A VGND VGND VPWR VPWR _0583_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1204_ _1211_/CLK _1204_/D VGND VGND VPWR VPWR _1204_/Q sky130_fd_sc_hd__dfxtp_1
X_1066_ _1195_/CLK _1066_/D VGND VGND VPWR VPWR _1066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1135_ _1195_/CLK _1135_/D VGND VGND VPWR VPWR _1135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0919_ _0926_/A VGND VGND VPWR VPWR _0919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0635_ _1173_/Q VGND VGND VPWR VPWR _0635_/Y sky130_fd_sc_hd__inv_2
X_0704_ _0798_/A VGND VGND VPWR VPWR _0704_/X sky130_fd_sc_hd__clkbuf_2
X_0566_ _1085_/Q VGND VGND VPWR VPWR _0566_/Y sky130_fd_sc_hd__inv_2
X_1049_ _1216_/CLK _1049_/D VGND VGND VPWR VPWR _1049_/Q sky130_fd_sc_hd__dfxtp_1
X_1118_ _1174_/CLK _1118_/D VGND VGND VPWR VPWR _1118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0618_ _1175_/Q VGND VGND VPWR VPWR _0618_/Y sky130_fd_sc_hd__inv_2
X_0549_ _0537_/X _1216_/Q _0511_/X _0548_/Y VGND VGND VPWR VPWR _1216_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0952_ _1089_/Q _0947_/X input44/X _0950_/X VGND VGND VPWR VPWR _1089_/D sky130_fd_sc_hd__a22o_1
Xoutput115 _1085_/Q VGND VGND VPWR VPWR o_cacheable_area[26] sky130_fd_sc_hd__clkbuf_2
Xoutput148 _1214_/Q VGND VGND VPWR VPWR o_copro_read_data[27] sky130_fd_sc_hd__clkbuf_2
Xoutput126 _1066_/Q VGND VGND VPWR VPWR o_cacheable_area[7] sky130_fd_sc_hd__clkbuf_2
Xoutput137 _1204_/Q VGND VGND VPWR VPWR o_copro_read_data[17] sky130_fd_sc_hd__clkbuf_2
Xoutput159 _1195_/Q VGND VGND VPWR VPWR o_copro_read_data[8] sky130_fd_sc_hd__clkbuf_2
X_0883_ _1131_/Q _0878_/X input51/X _0879_/X VGND VGND VPWR VPWR _1131_/D sky130_fd_sc_hd__a22o_1
Xoutput104 _1075_/Q VGND VGND VPWR VPWR o_cacheable_area[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput17 i_copro_opcode2[1] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_1
Xinput28 i_copro_write_data[16] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_2
Xinput39 i_copro_write_data[26] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1151_ _1215_/CLK _1151_/D VGND VGND VPWR VPWR _1151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1082_ _1180_/CLK _1082_/D VGND VGND VPWR VPWR _1082_/Q sky130_fd_sc_hd__dfxtp_2
X_0866_ _1144_/Q _0864_/X input34/X _0865_/X VGND VGND VPWR VPWR _1144_/D sky130_fd_sc_hd__a22o_1
X_0935_ _1097_/Q _0933_/X input83/X _0934_/X VGND VGND VPWR VPWR _1097_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0797_ _0797_/A VGND VGND VPWR VPWR _0944_/C sky130_fd_sc_hd__inv_2
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0720_ _1162_/Q VGND VGND VPWR VPWR _0720_/Y sky130_fd_sc_hd__inv_2
X_0651_ _0649_/Y _0594_/X _0650_/Y _0610_/X VGND VGND VPWR VPWR _0651_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0582_ _1147_/Q VGND VGND VPWR VPWR _0582_/Y sky130_fd_sc_hd__inv_2
X_1134_ _1166_/CLK _1134_/D VGND VGND VPWR VPWR _1134_/Q sky130_fd_sc_hd__dfxtp_1
X_1203_ _1211_/CLK _1203_/D VGND VGND VPWR VPWR _1203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1065_ _1187_/CLK _1065_/D VGND VGND VPWR VPWR _1065_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0918_ _1108_/Q _0912_/X input63/X _0913_/X VGND VGND VPWR VPWR _1108_/D sky130_fd_sc_hd__a22o_1
X_0849_ _0885_/A VGND VGND VPWR VPWR _0886_/A sky130_fd_sc_hd__inv_2
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0703_ _0663_/X _1197_/Q _0695_/X _0702_/Y VGND VGND VPWR VPWR _1197_/D sky130_fd_sc_hd__a22o_1
X_0565_ _1181_/Q VGND VGND VPWR VPWR _0565_/Y sky130_fd_sc_hd__inv_2
X_0634_ _1077_/Q VGND VGND VPWR VPWR _0634_/Y sky130_fd_sc_hd__inv_2
X_1117_ _1181_/CLK _1117_/D VGND VGND VPWR VPWR _1117_/Q sky130_fd_sc_hd__dfxtp_1
X_1048_ _1216_/CLK _1048_/D VGND VGND VPWR VPWR _1048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0617_ _0723_/A VGND VGND VPWR VPWR _0617_/X sky130_fd_sc_hd__clkbuf_2
X_0548_ _0538_/Y _0518_/X _0539_/Y _0541_/X _0547_/X VGND VGND VPWR VPWR _0548_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0882_ _1132_/Q _0878_/X input52/X _0879_/X VGND VGND VPWR VPWR _1132_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0951_ _1090_/Q _0947_/X input45/X _0950_/X VGND VGND VPWR VPWR _1090_/D sky130_fd_sc_hd__a22o_1
Xoutput149 _1215_/Q VGND VGND VPWR VPWR o_copro_read_data[28] sky130_fd_sc_hd__clkbuf_2
Xoutput127 _1067_/Q VGND VGND VPWR VPWR o_cacheable_area[8] sky130_fd_sc_hd__clkbuf_2
Xoutput138 _1205_/Q VGND VGND VPWR VPWR o_copro_read_data[18] sky130_fd_sc_hd__clkbuf_2
Xoutput116 _1086_/Q VGND VGND VPWR VPWR o_cacheable_area[27] sky130_fd_sc_hd__clkbuf_2
Xoutput105 _1076_/Q VGND VGND VPWR VPWR o_cacheable_area[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 i_copro_opcode2[2] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__buf_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput29 i_copro_write_data[17] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_2
X_1150_ _1215_/CLK _1150_/D VGND VGND VPWR VPWR _1150_/Q sky130_fd_sc_hd__dfxtp_1
X_1081_ _1181_/CLK _1081_/D VGND VGND VPWR VPWR _1081_/Q sky130_fd_sc_hd__dfxtp_2
X_0934_ _1001_/A VGND VGND VPWR VPWR _0934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0865_ _0865_/A VGND VGND VPWR VPWR _0865_/X sky130_fd_sc_hd__clkbuf_2
X_0796_ _0749_/X _1187_/Q _0614_/A _0795_/Y VGND VGND VPWR VPWR _1187_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0650_ _1139_/Q VGND VGND VPWR VPWR _0650_/Y sky130_fd_sc_hd__inv_2
X_0581_ _0625_/A VGND VGND VPWR VPWR _0581_/X sky130_fd_sc_hd__clkbuf_2
X_1133_ _1166_/CLK _1133_/D VGND VGND VPWR VPWR _1133_/Q sky130_fd_sc_hd__dfxtp_1
X_1202_ _1206_/CLK _1202_/D VGND VGND VPWR VPWR _1202_/Q sky130_fd_sc_hd__dfxtp_1
X_1064_ _1209_/CLK _1064_/D VGND VGND VPWR VPWR _1064_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0917_ _1109_/Q _0912_/X input64/X _0913_/X VGND VGND VPWR VPWR _1109_/D sky130_fd_sc_hd__a22o_1
X_0848_ _0864_/A VGND VGND VPWR VPWR _0848_/X sky130_fd_sc_hd__clkbuf_2
X_0779_ _1124_/Q VGND VGND VPWR VPWR _0779_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0702_ _0696_/Y _0697_/X _0698_/Y _0666_/X _0701_/X VGND VGND VPWR VPWR _0702_/Y
+ sky130_fd_sc_hd__o221ai_2
X_0633_ _1141_/Q VGND VGND VPWR VPWR _0633_/Y sky130_fd_sc_hd__inv_2
X_0564_ _0537_/X _1214_/Q _0511_/X _0563_/Y VGND VGND VPWR VPWR _1214_/D sky130_fd_sc_hd__a22o_1
X_1047_ _1056_/Q VGND VGND VPWR VPWR _1047_/X sky130_fd_sc_hd__buf_2
X_1116_ _1181_/CLK _1116_/D VGND VGND VPWR VPWR _1116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0616_ _1079_/Q VGND VGND VPWR VPWR _0616_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0547_ _0542_/Y _0544_/X _0545_/Y _0583_/A VGND VGND VPWR VPWR _0547_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0881_ _1133_/Q _0878_/X input22/X _0879_/X VGND VGND VPWR VPWR _1133_/D sky130_fd_sc_hd__a22o_1
X_0950_ _0964_/A VGND VGND VPWR VPWR _0950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput128 _1068_/Q VGND VGND VPWR VPWR o_cacheable_area[9] sky130_fd_sc_hd__clkbuf_2
Xoutput117 _1087_/Q VGND VGND VPWR VPWR o_cacheable_area[28] sky130_fd_sc_hd__clkbuf_2
Xoutput106 _1077_/Q VGND VGND VPWR VPWR o_cacheable_area[18] sky130_fd_sc_hd__clkbuf_2
Xoutput139 _1206_/Q VGND VGND VPWR VPWR o_copro_read_data[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 i_copro_operation[0] VGND VGND VPWR VPWR _0944_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ _1211_/CLK _1080_/D VGND VGND VPWR VPWR _1080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0933_ _1000_/A VGND VGND VPWR VPWR _0933_/X sky130_fd_sc_hd__clkbuf_2
X_0795_ _0787_/Y _0541_/A _0788_/Y _0583_/A _0794_/X VGND VGND VPWR VPWR _0795_/Y
+ sky130_fd_sc_hd__o221ai_1
X_0864_ _0864_/A VGND VGND VPWR VPWR _0864_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1201_ _1206_/CLK _1201_/D VGND VGND VPWR VPWR _1201_/Q sky130_fd_sc_hd__dfxtp_1
X_0580_ _0537_/X _1212_/Q _0572_/X _0579_/Y VGND VGND VPWR VPWR _1212_/D sky130_fd_sc_hd__a22o_1
X_1132_ _1166_/CLK _1132_/D VGND VGND VPWR VPWR _1132_/Q sky130_fd_sc_hd__dfxtp_1
X_1063_ _1209_/CLK _1063_/D VGND VGND VPWR VPWR _1063_/Q sky130_fd_sc_hd__dfxtp_2
X_0916_ _1110_/Q _0912_/X input65/X _0913_/X VGND VGND VPWR VPWR _1110_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0847_ _0885_/A VGND VGND VPWR VPWR _0864_/A sky130_fd_sc_hd__clkbuf_2
X_0778_ _1060_/Q VGND VGND VPWR VPWR _0778_/Y sky130_fd_sc_hd__inv_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0701_ _0699_/Y _0668_/X _0700_/Y _0677_/X VGND VGND VPWR VPWR _0701_/X sky130_fd_sc_hd__o22a_1
X_0632_ _0625_/X _1206_/Q _0614_/X _0631_/Y VGND VGND VPWR VPWR _1206_/D sky130_fd_sc_hd__a22o_1
X_0563_ _0558_/Y _0518_/X _0559_/Y _0541_/X _0562_/X VGND VGND VPWR VPWR _0563_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1046_ _1090_/Q VGND VGND VPWR VPWR _1046_/X sky130_fd_sc_hd__buf_2
X_1115_ _1181_/CLK _1115_/D VGND VGND VPWR VPWR _1115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0615_ _1143_/Q VGND VGND VPWR VPWR _0615_/Y sky130_fd_sc_hd__inv_2
X_0546_ _0846_/D VGND VGND VPWR VPWR _0583_/A sky130_fd_sc_hd__buf_2
X_1029_ _1073_/Q VGND VGND VPWR VPWR _1029_/X sky130_fd_sc_hd__buf_2
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0529_ _0993_/A input6/X input8/X _0726_/B VGND VGND VPWR VPWR _0846_/D sky130_fd_sc_hd__or4_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput107 _1078_/Q VGND VGND VPWR VPWR o_cacheable_area[19] sky130_fd_sc_hd__clkbuf_2
X_0880_ _1134_/Q _0878_/X input23/X _0879_/X VGND VGND VPWR VPWR _1134_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput118 _1088_/Q VGND VGND VPWR VPWR o_cacheable_area[29] sky130_fd_sc_hd__clkbuf_2
Xoutput129 _1187_/Q VGND VGND VPWR VPWR o_copro_read_data[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0932_ _1098_/Q _0926_/X input84/X _0927_/X VGND VGND VPWR VPWR _1098_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0863_ _1145_/Q _0857_/X input35/X _0858_/X VGND VGND VPWR VPWR _1145_/D sky130_fd_sc_hd__a22o_1
X_0794_ _0789_/Y _0602_/A _0790_/Y _0770_/X _0793_/X VGND VGND VPWR VPWR _0794_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1200_ _1200_/CLK _1200_/D VGND VGND VPWR VPWR _1200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1131_ _1166_/CLK _1131_/D VGND VGND VPWR VPWR _1131_/Q sky130_fd_sc_hd__dfxtp_1
X_1062_ _1209_/CLK _1062_/D VGND VGND VPWR VPWR _1062_/Q sky130_fd_sc_hd__dfxtp_2
X_0915_ _1111_/Q _0912_/X input67/X _0913_/X VGND VGND VPWR VPWR _1111_/D sky130_fd_sc_hd__a22o_1
X_0846_ _0944_/A _0944_/B _0944_/C _0846_/D VGND VGND VPWR VPWR _0885_/A sky130_fd_sc_hd__or4_4
X_0777_ _1049_/Q VGND VGND VPWR VPWR _0777_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0700_ _1133_/Q VGND VGND VPWR VPWR _0700_/Y sky130_fd_sc_hd__inv_2
X_0631_ _0626_/Y _0574_/X _0627_/Y _0592_/X _0630_/X VGND VGND VPWR VPWR _0631_/Y
+ sky130_fd_sc_hd__o221ai_4
X_0562_ _0560_/Y _0544_/X _0561_/Y _0554_/X VGND VGND VPWR VPWR _0562_/X sky130_fd_sc_hd__o22a_1
X_1114_ _1181_/CLK _1114_/D VGND VGND VPWR VPWR _1114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1045_ _1089_/Q VGND VGND VPWR VPWR _1045_/X sky130_fd_sc_hd__buf_2
X_0829_ _1167_/Q _0823_/X input24/X _0824_/X VGND VGND VPWR VPWR _1167_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_i_clk clkbuf_3_6_0_i_clk/X VGND VGND VPWR VPWR _1170_/CLK sky130_fd_sc_hd__clkbuf_1
X_0545_ _1152_/Q VGND VGND VPWR VPWR _0545_/Y sky130_fd_sc_hd__inv_2
X_0614_ _0614_/A VGND VGND VPWR VPWR _0614_/X sky130_fd_sc_hd__clkbuf_2
X_1028_ _1072_/Q VGND VGND VPWR VPWR _1028_/X sky130_fd_sc_hd__buf_2
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0528_ _1153_/Q VGND VGND VPWR VPWR _0528_/Y sky130_fd_sc_hd__inv_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput108 _1060_/Q VGND VGND VPWR VPWR o_cacheable_area[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput119 _1061_/Q VGND VGND VPWR VPWR o_cacheable_area[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0931_ _1099_/Q _0926_/X input85/X _0927_/X VGND VGND VPWR VPWR _1099_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0862_ _1146_/Q _0857_/X input36/X _0858_/X VGND VGND VPWR VPWR _1146_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0793_ _0791_/Y _0736_/A _0792_/Y _0798_/D VGND VGND VPWR VPWR _0793_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1130_ _1195_/CLK _1130_/D VGND VGND VPWR VPWR _1130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1061_ _1216_/CLK _1061_/D VGND VGND VPWR VPWR _1061_/Q sky130_fd_sc_hd__dfxtp_2
X_0914_ _1112_/Q _0912_/X input68/X _0913_/X VGND VGND VPWR VPWR _1112_/D sky130_fd_sc_hd__a22o_1
X_0845_ _1155_/Q _0816_/A input21/X _0817_/A VGND VGND VPWR VPWR _1155_/D sky130_fd_sc_hd__a22o_1
X_0776_ _0749_/X _1189_/Q _0740_/X _0775_/Y VGND VGND VPWR VPWR _1189_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0630_ _0628_/Y _0594_/X _0629_/Y _0610_/X VGND VGND VPWR VPWR _0630_/X sky130_fd_sc_hd__o22a_1
X_0561_ _1150_/Q VGND VGND VPWR VPWR _0561_/Y sky130_fd_sc_hd__inv_2
X_1044_ _1088_/Q VGND VGND VPWR VPWR _1044_/X sky130_fd_sc_hd__buf_2
X_1113_ _1181_/CLK _1113_/D VGND VGND VPWR VPWR _1113_/Q sky130_fd_sc_hd__dfxtp_1
X_0828_ _1168_/Q _0823_/X input25/X _0824_/X VGND VGND VPWR VPWR _1168_/D sky130_fd_sc_hd__a22o_1
X_0759_ _1126_/Q VGND VGND VPWR VPWR _0759_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0613_ _0581_/X _1208_/Q _0572_/X _0612_/Y VGND VGND VPWR VPWR _1208_/D sky130_fd_sc_hd__a22o_1
X_0544_ _0668_/A VGND VGND VPWR VPWR _0544_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1027_ _1071_/Q VGND VGND VPWR VPWR _1027_/X sky130_fd_sc_hd__buf_2
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0527_ _0723_/A VGND VGND VPWR VPWR _0666_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput109 _1079_/Q VGND VGND VPWR VPWR o_cacheable_area[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0930_ _1100_/Q _0926_/X input86/X _0927_/X VGND VGND VPWR VPWR _1100_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0792_ _1155_/Q VGND VGND VPWR VPWR _0792_/Y sky130_fd_sc_hd__inv_2
X_0861_ _1147_/Q _0857_/X input37/X _0858_/X VGND VGND VPWR VPWR _1147_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_3_7_0_i_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1060_ _1170_/CLK _1060_/D VGND VGND VPWR VPWR _1060_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0913_ _0927_/A VGND VGND VPWR VPWR _0913_/X sky130_fd_sc_hd__clkbuf_2
X_0844_ _1156_/Q _0816_/A input32/X _0817_/A VGND VGND VPWR VPWR _1156_/D sky130_fd_sc_hd__a22o_1
X_0775_ _0766_/Y _0736_/A _0767_/Y _0541_/A _0774_/X VGND VGND VPWR VPWR _0775_/Y
+ sky130_fd_sc_hd__o221ai_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1189_ _1210_/CLK _1189_/D VGND VGND VPWR VPWR _1189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0560_ _1118_/Q VGND VGND VPWR VPWR _0560_/Y sky130_fd_sc_hd__inv_2
X_1112_ _1166_/CLK _1112_/D VGND VGND VPWR VPWR _1112_/Q sky130_fd_sc_hd__dfxtp_1
X_1043_ _1087_/Q VGND VGND VPWR VPWR _1043_/X sky130_fd_sc_hd__buf_2
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0827_ _1169_/Q _0823_/X input26/X _0824_/X VGND VGND VPWR VPWR _1169_/D sky130_fd_sc_hd__a22o_1
X_0758_ _1158_/Q VGND VGND VPWR VPWR _0758_/Y sky130_fd_sc_hd__inv_2
X_0689_ _1070_/Q VGND VGND VPWR VPWR _0689_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0612_ _0606_/Y _0574_/X _0607_/Y _0592_/X _0611_/X VGND VGND VPWR VPWR _0612_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0543_ _0725_/A VGND VGND VPWR VPWR _0668_/A sky130_fd_sc_hd__clkbuf_2
X_1026_ _1070_/Q VGND VGND VPWR VPWR _1026_/X sky130_fd_sc_hd__buf_2
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_i_clk clkbuf_4_7_0_i_clk/A VGND VGND VPWR VPWR _1211_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0526_ _1007_/A _0993_/B _0944_/D VGND VGND VPWR VPWR _0723_/A sky130_fd_sc_hd__or3_4
XANTENNA_0 input21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1090_/Q VGND VGND VPWR VPWR _1009_/Y sky130_fd_sc_hd__inv_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0509_ _0944_/A VGND VGND VPWR VPWR _0894_/A sky130_fd_sc_hd__inv_2
XFILLER_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_i_clk clkbuf_0_i_clk/X VGND VGND VPWR VPWR clkbuf_4_7_0_i_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0791_ _1048_/Q VGND VGND VPWR VPWR _0791_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0860_ _1148_/Q _0857_/X input38/X _0858_/X VGND VGND VPWR VPWR _1148_/D sky130_fd_sc_hd__a22o_1
X_0989_ _1062_/Q _0984_/X input46/X _0985_/X VGND VGND VPWR VPWR _1062_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0912_ _0926_/A VGND VGND VPWR VPWR _0912_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0843_ _1157_/Q _0837_/X input43/X _0838_/X VGND VGND VPWR VPWR _1157_/D sky130_fd_sc_hd__a22o_1
X_0774_ _0768_/Y _0706_/A _0769_/Y _0770_/X _0773_/X VGND VGND VPWR VPWR _0774_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ _1210_/CLK _1188_/D VGND VGND VPWR VPWR _1188_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1111_ _1166_/CLK _1111_/D VGND VGND VPWR VPWR _1111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1042_ _1086_/Q VGND VGND VPWR VPWR _1042_/X sky130_fd_sc_hd__buf_2
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0688_ _1166_/Q VGND VGND VPWR VPWR _0688_/Y sky130_fd_sc_hd__inv_2
X_0826_ _1170_/Q _0823_/X input27/X _0824_/X VGND VGND VPWR VPWR _1170_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_4_2_0_i_clk clkbuf_4_3_0_i_clk/A VGND VGND VPWR VPWR _1215_/CLK sky130_fd_sc_hd__clkbuf_1
X_0757_ _0749_/X _1191_/Q _0740_/X _0756_/Y VGND VGND VPWR VPWR _1191_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0611_ _0608_/Y _0594_/X _0609_/Y _0610_/X VGND VGND VPWR VPWR _0611_/X sky130_fd_sc_hd__o22a_1
X_0542_ _1120_/Q VGND VGND VPWR VPWR _0542_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1025_ _1069_/Q VGND VGND VPWR VPWR _1025_/X sky130_fd_sc_hd__buf_2
X_0809_ _0816_/A VGND VGND VPWR VPWR _0809_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0525_ _0726_/D VGND VGND VPWR VPWR _0993_/B sky130_fd_sc_hd__buf_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1008_ _1186_/Q VGND VGND VPWR VPWR _1008_/Y sky130_fd_sc_hd__inv_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0508_ _0798_/A VGND VGND VPWR VPWR _0625_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0790_ _1056_/Q VGND VGND VPWR VPWR _0790_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0988_ _1063_/Q _0984_/X input47/X _0985_/X VGND VGND VPWR VPWR _1063_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0911_ _1113_/Q _0905_/X input69/X _0906_/X VGND VGND VPWR VPWR _1113_/D sky130_fd_sc_hd__a22o_1
X_0842_ _1158_/Q _0837_/X input46/X _0838_/X VGND VGND VPWR VPWR _1158_/D sky130_fd_sc_hd__a22o_1
X_0773_ _0771_/Y _0668_/A _0772_/Y _0697_/A VGND VGND VPWR VPWR _0773_/X sky130_fd_sc_hd__o22a_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1187_ _1187_/CLK _1187_/D VGND VGND VPWR VPWR _1187_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1110_ _1176_/CLK _1110_/D VGND VGND VPWR VPWR _1110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1041_ _1085_/Q VGND VGND VPWR VPWR _1041_/X sky130_fd_sc_hd__buf_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0825_ _1171_/Q _0823_/X input28/X _0824_/X VGND VGND VPWR VPWR _1171_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0687_ _0663_/X _1199_/Q _0654_/X _0686_/Y VGND VGND VPWR VPWR _1199_/D sky130_fd_sc_hd__a22o_1
X_0756_ _0750_/Y _0697_/X _0751_/Y _0583_/A _0755_/X VGND VGND VPWR VPWR _0756_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0610_ _0846_/D VGND VGND VPWR VPWR _0610_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0541_ _0541_/A VGND VGND VPWR VPWR _0541_/X sky130_fd_sc_hd__buf_2
X_1024_ _1068_/Q VGND VGND VPWR VPWR _1024_/X sky130_fd_sc_hd__buf_2
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0808_ _1182_/Q _0800_/X input40/X _0803_/X VGND VGND VPWR VPWR _1182_/D sky130_fd_sc_hd__a22o_1
X_0739_ _0704_/X _1193_/Q _0695_/X _0738_/Y VGND VGND VPWR VPWR _1193_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0524_ input6/X VGND VGND VPWR VPWR _0726_/D sky130_fd_sc_hd__inv_2
X_1007_ _1007_/A input6/X _1007_/C VGND VGND VPWR VPWR _1007_/Y sky130_fd_sc_hd__nor3_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0507_ _0944_/A VGND VGND VPWR VPWR _0798_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0987_ _1064_/Q _0984_/X input48/X _0985_/X VGND VGND VPWR VPWR _1064_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0910_ _1114_/Q _0905_/X input70/X _0906_/X VGND VGND VPWR VPWR _1114_/D sky130_fd_sc_hd__a22o_1
X_0841_ _1159_/Q _0837_/X input47/X _0838_/X VGND VGND VPWR VPWR _1159_/D sky130_fd_sc_hd__a22o_1
X_0772_ _1157_/Q VGND VGND VPWR VPWR _0772_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1186_ _1218_/CLK _1186_/D VGND VGND VPWR VPWR _1186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1040_ _1084_/Q VGND VGND VPWR VPWR _1040_/X sky130_fd_sc_hd__buf_2
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0824_ _0838_/A VGND VGND VPWR VPWR _0824_/X sky130_fd_sc_hd__buf_1
X_0755_ _0752_/Y _0723_/X _0753_/Y _0725_/X _0754_/X VGND VGND VPWR VPWR _0755_/X
+ sky130_fd_sc_hd__o221a_1
X_0686_ _0681_/Y _0656_/X _0682_/Y _0666_/X _0685_/X VGND VGND VPWR VPWR _0686_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1169_ _1206_/CLK _1169_/D VGND VGND VPWR VPWR _1169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0540_ _0723_/A VGND VGND VPWR VPWR _0541_/A sky130_fd_sc_hd__buf_2
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1023_ _1067_/Q VGND VGND VPWR VPWR _1023_/X sky130_fd_sc_hd__buf_2
X_0807_ _1183_/Q _0800_/X input41/X _0803_/X VGND VGND VPWR VPWR _1183_/D sky130_fd_sc_hd__a22o_1
X_0738_ _0732_/Y _0697_/X _0733_/Y _0706_/X _0737_/X VGND VGND VPWR VPWR _0738_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0669_ _1137_/Q VGND VGND VPWR VPWR _0669_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0523_ _1089_/Q VGND VGND VPWR VPWR _0523_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1006_ _1048_/Q _1000_/X input87/X _1001_/X VGND VGND VPWR VPWR _1048_/D sky130_fd_sc_hd__a22o_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput95 _1056_/Q VGND VGND VPWR VPWR o_cache_enable sky130_fd_sc_hd__clkbuf_2
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0986_ _1065_/Q _0984_/X input49/X _0985_/X VGND VGND VPWR VPWR _1065_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0771_ _1093_/Q VGND VGND VPWR VPWR _0771_/Y sky130_fd_sc_hd__inv_2
X_0840_ _1160_/Q _0837_/X input48/X _0838_/X VGND VGND VPWR VPWR _1160_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1185_ _1218_/CLK _1185_/D VGND VGND VPWR VPWR _1185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0969_ _1076_/Q _0963_/X input29/X _0964_/X VGND VGND VPWR VPWR _1076_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0685_ _0683_/Y _0668_/X _0684_/Y _0677_/X VGND VGND VPWR VPWR _0685_/X sky130_fd_sc_hd__o22a_1
X_0823_ _0837_/A VGND VGND VPWR VPWR _0823_/X sky130_fd_sc_hd__clkbuf_2
X_0754_ _0762_/A _1052_/Q VGND VGND VPWR VPWR _0754_/X sky130_fd_sc_hd__or2b_1
X_1099_ _1176_/CLK _1099_/D VGND VGND VPWR VPWR _1099_/Q sky130_fd_sc_hd__dfxtp_1
X_1168_ _1206_/CLK _1168_/D VGND VGND VPWR VPWR _1168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1022_ _1066_/Q VGND VGND VPWR VPWR _1022_/X sky130_fd_sc_hd__buf_2
X_0668_ _0668_/A VGND VGND VPWR VPWR _0668_/X sky130_fd_sc_hd__clkbuf_2
X_0806_ _1184_/Q _0800_/X input42/X _0803_/X VGND VGND VPWR VPWR _1184_/D sky130_fd_sc_hd__a22o_1
X_0737_ _0734_/Y _0723_/X _0735_/Y _0725_/X _0736_/X VGND VGND VPWR VPWR _0737_/X
+ sky130_fd_sc_hd__o221a_1
X_0599_ _1145_/Q VGND VGND VPWR VPWR _0599_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0522_ _0522_/A VGND VGND VPWR VPWR _0522_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ _1049_/Q _1000_/X input88/X _1001_/X VGND VGND VPWR VPWR _1049_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput96 _1007_/Y VGND VGND VPWR VPWR o_cache_flush sky130_fd_sc_hd__clkbuf_2
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

