magic
tech sky130A
magscale 1 2
timestamp 1618216021
<< checkpaint >>
rect -3932 -3932 33512 35656
<< locali >>
rect 9505 26775 9539 27081
rect 10333 20927 10367 21097
rect 21741 20791 21775 21029
rect 5917 18615 5951 18853
rect 8953 18751 8987 18853
rect 14197 18615 14231 18921
rect 14565 15895 14599 16065
rect 3433 13855 3467 13957
rect 20361 7871 20395 8041
rect 20361 7735 20395 7837
<< viali >>
rect 4445 29257 4479 29291
rect 7113 29257 7147 29291
rect 7849 29257 7883 29291
rect 10793 29257 10827 29291
rect 13369 29257 13403 29291
rect 16589 29257 16623 29291
rect 18797 29257 18831 29291
rect 20913 29257 20947 29291
rect 21833 29257 21867 29291
rect 23857 29257 23891 29291
rect 24593 29257 24627 29291
rect 2697 29189 2731 29223
rect 5825 29189 5859 29223
rect 8677 29189 8711 29223
rect 15945 29189 15979 29223
rect 23213 29189 23247 29223
rect 25881 29189 25915 29223
rect 27353 29121 27387 29155
rect 1869 29053 1903 29087
rect 2513 29053 2547 29087
rect 7021 29053 7055 29087
rect 9965 29053 9999 29087
rect 10149 29053 10183 29087
rect 12541 29053 12575 29087
rect 13277 29053 13311 29087
rect 15025 29053 15059 29087
rect 15209 29053 15243 29087
rect 16405 29053 16439 29087
rect 17601 29053 17635 29087
rect 17785 29053 17819 29087
rect 18015 29053 18049 29087
rect 18705 29053 18739 29087
rect 21741 29053 21775 29087
rect 23029 29053 23063 29087
rect 24501 29053 24535 29087
rect 26433 29053 26467 29087
rect 27169 29053 27203 29087
rect 2053 28985 2087 29019
rect 4353 28985 4387 29019
rect 5641 28985 5675 29019
rect 7757 28985 7791 29019
rect 8493 28985 8527 29019
rect 10701 28985 10735 29019
rect 12725 28985 12759 29019
rect 15761 28985 15795 29019
rect 17873 28985 17907 29019
rect 20821 28985 20855 29019
rect 23765 28985 23799 29019
rect 25697 28985 25731 29019
rect 26617 28985 26651 29019
rect 18153 28917 18187 28951
rect 1961 28713 1995 28747
rect 3065 28713 3099 28747
rect 16129 28713 16163 28747
rect 7481 28645 7515 28679
rect 24317 28645 24351 28679
rect 25789 28645 25823 28679
rect 1869 28577 1903 28611
rect 2973 28577 3007 28611
rect 4261 28577 4295 28611
rect 5089 28577 5123 28611
rect 6193 28577 6227 28611
rect 7297 28577 7331 28611
rect 7573 28577 7607 28611
rect 7711 28577 7745 28611
rect 8309 28577 8343 28611
rect 9505 28577 9539 28611
rect 10508 28577 10542 28611
rect 12081 28577 12115 28611
rect 12909 28577 12943 28611
rect 13369 28577 13403 28611
rect 15016 28577 15050 28611
rect 16589 28577 16623 28611
rect 17776 28577 17810 28611
rect 20085 28577 20119 28611
rect 20821 28577 20855 28611
rect 21557 28577 21591 28611
rect 22293 28577 22327 28611
rect 23397 28577 23431 28611
rect 24133 28577 24167 28611
rect 25605 28577 25639 28611
rect 26341 28577 26375 28611
rect 26985 28577 27019 28611
rect 10241 28509 10275 28543
rect 14749 28509 14783 28543
rect 17509 28509 17543 28543
rect 5273 28441 5307 28475
rect 22477 28441 22511 28475
rect 4445 28373 4479 28407
rect 7849 28373 7883 28407
rect 8493 28373 8527 28407
rect 11621 28373 11655 28407
rect 12725 28373 12759 28407
rect 18889 28373 18923 28407
rect 23581 28373 23615 28407
rect 26433 28373 26467 28407
rect 2329 28169 2363 28203
rect 2973 28101 3007 28135
rect 18889 28101 18923 28135
rect 1409 27965 1443 27999
rect 2145 27965 2179 27999
rect 2789 27965 2823 27999
rect 3617 27965 3651 27999
rect 6837 27965 6871 27999
rect 7104 27965 7138 27999
rect 8677 27965 8711 27999
rect 10517 27965 10551 27999
rect 12081 27965 12115 27999
rect 13921 27965 13955 27999
rect 14381 27965 14415 27999
rect 17509 27965 17543 27999
rect 17776 27965 17810 27999
rect 19349 27965 19383 27999
rect 20269 27965 20303 27999
rect 20453 27965 20487 27999
rect 20545 27965 20579 27999
rect 20637 27965 20671 27999
rect 21281 27965 21315 27999
rect 22569 27965 22603 27999
rect 23949 27965 23983 27999
rect 24593 27965 24627 27999
rect 25329 27965 25363 27999
rect 25973 27965 26007 27999
rect 26709 27965 26743 27999
rect 8922 27897 8956 27931
rect 14648 27897 14682 27931
rect 3433 27829 3467 27863
rect 8217 27829 8251 27863
rect 10057 27829 10091 27863
rect 12265 27829 12299 27863
rect 13737 27829 13771 27863
rect 15761 27829 15795 27863
rect 20821 27829 20855 27863
rect 22753 27829 22787 27863
rect 24133 27829 24167 27863
rect 10701 27625 10735 27659
rect 15301 27625 15335 27659
rect 16313 27625 16347 27659
rect 18061 27625 18095 27659
rect 10333 27557 10367 27591
rect 15025 27557 15059 27591
rect 15945 27557 15979 27591
rect 17693 27557 17727 27591
rect 17785 27557 17819 27591
rect 20628 27557 20662 27591
rect 25789 27557 25823 27591
rect 26525 27557 26559 27591
rect 1961 27489 1995 27523
rect 6644 27489 6678 27523
rect 8217 27489 8251 27523
rect 9505 27489 9539 27523
rect 10149 27489 10183 27523
rect 10425 27489 10459 27523
rect 10517 27489 10551 27523
rect 12164 27489 12198 27523
rect 14749 27489 14783 27523
rect 14933 27489 14967 27523
rect 15117 27489 15151 27523
rect 15761 27489 15795 27523
rect 16037 27489 16071 27523
rect 16129 27489 16163 27523
rect 16773 27489 16807 27523
rect 17509 27489 17543 27523
rect 17877 27489 17911 27523
rect 18521 27489 18555 27523
rect 25605 27489 25639 27523
rect 26341 27489 26375 27523
rect 26985 27489 27019 27523
rect 6377 27421 6411 27455
rect 11897 27421 11931 27455
rect 20361 27421 20395 27455
rect 21741 27353 21775 27387
rect 1777 27285 1811 27319
rect 7757 27285 7791 27319
rect 9597 27285 9631 27319
rect 13277 27285 13311 27319
rect 16957 27285 16991 27319
rect 18705 27285 18739 27319
rect 7665 27081 7699 27115
rect 8677 27081 8711 27115
rect 9505 27081 9539 27115
rect 2145 26877 2179 26911
rect 7113 26877 7147 26911
rect 7389 26877 7423 26911
rect 7481 26877 7515 26911
rect 8125 26877 8159 26911
rect 8493 26877 8527 26911
rect 7297 26809 7331 26843
rect 8309 26809 8343 26843
rect 8401 26809 8435 26843
rect 10609 27013 10643 27047
rect 26893 27013 26927 27047
rect 9597 26877 9631 26911
rect 9873 26877 9907 26911
rect 9965 26877 9999 26911
rect 10793 26877 10827 26911
rect 12081 26877 12115 26911
rect 13921 26877 13955 26911
rect 15025 26877 15059 26911
rect 15209 26877 15243 26911
rect 15393 26877 15427 26911
rect 16129 26877 16163 26911
rect 17325 26877 17359 26911
rect 17509 26877 17543 26911
rect 17693 26877 17727 26911
rect 18337 26877 18371 26911
rect 18981 26877 19015 26911
rect 21465 26877 21499 26911
rect 22845 26877 22879 26911
rect 23121 26877 23155 26911
rect 23213 26877 23247 26911
rect 9781 26809 9815 26843
rect 12348 26809 12382 26843
rect 15301 26809 15335 26843
rect 17601 26809 17635 26843
rect 23029 26809 23063 26843
rect 26709 26809 26743 26843
rect 9505 26741 9539 26775
rect 10149 26741 10183 26775
rect 13461 26741 13495 26775
rect 14013 26741 14047 26775
rect 15577 26741 15611 26775
rect 16221 26741 16255 26775
rect 17877 26741 17911 26775
rect 18429 26741 18463 26775
rect 19073 26741 19107 26775
rect 21557 26741 21591 26775
rect 23397 26741 23431 26775
rect 1961 26537 1995 26571
rect 16497 26537 16531 26571
rect 18521 26537 18555 26571
rect 22293 26537 22327 26571
rect 24317 26537 24351 26571
rect 9772 26469 9806 26503
rect 12072 26469 12106 26503
rect 15384 26469 15418 26503
rect 17408 26469 17442 26503
rect 23204 26469 23238 26503
rect 26801 26469 26835 26503
rect 27721 26469 27755 26503
rect 1869 26401 1903 26435
rect 11805 26401 11839 26435
rect 13645 26401 13679 26435
rect 15117 26401 15151 26435
rect 17141 26401 17175 26435
rect 20913 26401 20947 26435
rect 21180 26401 21214 26435
rect 27537 26401 27571 26435
rect 9505 26333 9539 26367
rect 22937 26333 22971 26367
rect 13737 26265 13771 26299
rect 26985 26265 27019 26299
rect 10885 26197 10919 26231
rect 13185 26197 13219 26231
rect 7113 25993 7147 26027
rect 7849 25993 7883 26027
rect 12633 25993 12667 26027
rect 21465 25993 21499 26027
rect 24225 25993 24259 26027
rect 14749 25925 14783 25959
rect 1685 25857 1719 25891
rect 14473 25857 14507 25891
rect 26893 25857 26927 25891
rect 1501 25789 1535 25823
rect 2145 25789 2179 25823
rect 2881 25789 2915 25823
rect 5273 25789 5307 25823
rect 5457 25789 5491 25823
rect 5641 25789 5675 25823
rect 6837 25789 6871 25823
rect 7757 25789 7791 25823
rect 9781 25789 9815 25823
rect 12081 25789 12115 25823
rect 12357 25789 12391 25823
rect 12449 25789 12483 25823
rect 13553 25789 13587 25823
rect 13829 25789 13863 25823
rect 14197 25789 14231 25823
rect 14749 25789 14783 25823
rect 15853 25789 15887 25823
rect 16037 25789 16071 25823
rect 16129 25789 16163 25823
rect 16221 25789 16255 25823
rect 17325 25789 17359 25823
rect 20913 25789 20947 25823
rect 21281 25789 21315 25823
rect 22845 25789 22879 25823
rect 24685 25789 24719 25823
rect 25053 25789 25087 25823
rect 26709 25789 26743 25823
rect 3148 25721 3182 25755
rect 5549 25721 5583 25755
rect 10048 25721 10082 25755
rect 12265 25721 12299 25755
rect 17570 25721 17604 25755
rect 21097 25721 21131 25755
rect 21189 25721 21223 25755
rect 23112 25721 23146 25755
rect 24869 25721 24903 25755
rect 24961 25721 24995 25755
rect 4261 25653 4295 25687
rect 5825 25653 5859 25687
rect 7297 25653 7331 25687
rect 11161 25653 11195 25687
rect 16405 25653 16439 25687
rect 18705 25653 18739 25687
rect 25237 25653 25271 25687
rect 3341 25449 3375 25483
rect 6561 25449 6595 25483
rect 11437 25449 11471 25483
rect 12817 25449 12851 25483
rect 13829 25449 13863 25483
rect 23397 25449 23431 25483
rect 26617 25449 26651 25483
rect 2973 25381 3007 25415
rect 3065 25381 3099 25415
rect 5448 25381 5482 25415
rect 11161 25381 11195 25415
rect 12449 25381 12483 25415
rect 12541 25381 12575 25415
rect 13553 25381 13587 25415
rect 15016 25381 15050 25415
rect 23121 25381 23155 25415
rect 25482 25381 25516 25415
rect 1409 25313 1443 25347
rect 2789 25313 2823 25347
rect 3157 25313 3191 25347
rect 4261 25313 4295 25347
rect 7113 25313 7147 25347
rect 7251 25313 7285 25347
rect 7389 25313 7423 25347
rect 7481 25313 7515 25347
rect 8125 25313 8159 25347
rect 9505 25313 9539 25347
rect 10149 25313 10183 25347
rect 10885 25313 10919 25347
rect 11069 25313 11103 25347
rect 11253 25313 11287 25347
rect 12265 25313 12299 25347
rect 12633 25313 12667 25347
rect 13277 25313 13311 25347
rect 13461 25313 13495 25347
rect 13645 25313 13679 25347
rect 14749 25313 14783 25347
rect 16681 25313 16715 25347
rect 17325 25313 17359 25347
rect 17785 25313 17819 25347
rect 18153 25313 18187 25347
rect 18337 25313 18371 25347
rect 18797 25313 18831 25347
rect 22845 25313 22879 25347
rect 23029 25313 23063 25347
rect 23213 25313 23247 25347
rect 27077 25313 27111 25347
rect 5181 25245 5215 25279
rect 16773 25245 16807 25279
rect 17509 25245 17543 25279
rect 25237 25245 25271 25279
rect 8585 25177 8619 25211
rect 17877 25177 17911 25211
rect 1593 25109 1627 25143
rect 4353 25109 4387 25143
rect 7665 25109 7699 25143
rect 8217 25109 8251 25143
rect 9597 25109 9631 25143
rect 10241 25109 10275 25143
rect 16129 25109 16163 25143
rect 18889 25109 18923 25143
rect 18889 24905 18923 24939
rect 5365 24837 5399 24871
rect 7205 24837 7239 24871
rect 13277 24837 13311 24871
rect 14473 24837 14507 24871
rect 18061 24837 18095 24871
rect 23581 24837 23615 24871
rect 7665 24769 7699 24803
rect 10333 24769 10367 24803
rect 10793 24769 10827 24803
rect 12725 24769 12759 24803
rect 14013 24769 14047 24803
rect 15577 24769 15611 24803
rect 16313 24769 16347 24803
rect 17509 24769 17543 24803
rect 2237 24701 2271 24735
rect 2605 24701 2639 24735
rect 3249 24701 3283 24735
rect 10057 24701 10091 24735
rect 10241 24701 10275 24735
rect 10425 24701 10459 24735
rect 10609 24701 10643 24735
rect 12081 24701 12115 24735
rect 12173 24701 12207 24735
rect 13001 24701 13035 24735
rect 13277 24701 13311 24735
rect 14197 24701 14231 24735
rect 14289 24701 14323 24735
rect 14565 24701 14599 24735
rect 15301 24701 15335 24735
rect 15393 24701 15427 24735
rect 15669 24701 15703 24735
rect 16221 24701 16255 24735
rect 17325 24701 17359 24735
rect 17785 24701 17819 24735
rect 18153 24701 18187 24735
rect 18337 24701 18371 24735
rect 18797 24701 18831 24735
rect 21189 24701 21223 24735
rect 23029 24701 23063 24735
rect 23213 24701 23247 24735
rect 23397 24701 23431 24735
rect 24041 24701 24075 24735
rect 26157 24701 26191 24735
rect 26525 24701 26559 24735
rect 1593 24633 1627 24667
rect 2421 24633 2455 24667
rect 2513 24633 2547 24667
rect 3516 24633 3550 24667
rect 5181 24633 5215 24667
rect 7021 24633 7055 24667
rect 7932 24633 7966 24667
rect 13553 24633 13587 24667
rect 15117 24633 15151 24667
rect 23305 24633 23339 24667
rect 24286 24633 24320 24667
rect 26341 24633 26375 24667
rect 26433 24633 26467 24667
rect 1685 24565 1719 24599
rect 2789 24565 2823 24599
rect 4629 24565 4663 24599
rect 9045 24565 9079 24599
rect 21281 24565 21315 24599
rect 25421 24565 25455 24599
rect 26709 24565 26743 24599
rect 3341 24361 3375 24395
rect 4813 24361 4847 24395
rect 8585 24361 8619 24395
rect 13185 24361 13219 24395
rect 15301 24361 15335 24395
rect 27445 24361 27479 24395
rect 2228 24293 2262 24327
rect 4537 24293 4571 24327
rect 5549 24293 5583 24327
rect 6368 24293 6402 24327
rect 8309 24293 8343 24327
rect 14933 24293 14967 24327
rect 15025 24293 15059 24327
rect 17509 24293 17543 24327
rect 22753 24293 22787 24327
rect 25513 24293 25547 24327
rect 26332 24293 26366 24327
rect 1961 24225 1995 24259
rect 4261 24225 4295 24259
rect 4445 24225 4479 24259
rect 4629 24225 4663 24259
rect 5365 24225 5399 24259
rect 8033 24225 8067 24259
rect 8217 24225 8251 24259
rect 8401 24225 8435 24259
rect 9873 24225 9907 24259
rect 10129 24225 10163 24259
rect 13093 24225 13127 24259
rect 14749 24225 14783 24259
rect 15117 24225 15151 24259
rect 15761 24225 15795 24259
rect 20545 24225 20579 24259
rect 21281 24225 21315 24259
rect 21741 24225 21775 24259
rect 22109 24225 22143 24259
rect 22293 24225 22327 24259
rect 22937 24225 22971 24259
rect 23029 24225 23063 24259
rect 23305 24225 23339 24259
rect 25421 24225 25455 24259
rect 6101 24157 6135 24191
rect 15853 24157 15887 24191
rect 20637 24157 20671 24191
rect 21465 24157 21499 24191
rect 26065 24157 26099 24191
rect 17693 24089 17727 24123
rect 22017 24089 22051 24123
rect 7481 24021 7515 24055
rect 11253 24021 11287 24055
rect 23213 24021 23247 24055
rect 5733 23817 5767 23851
rect 19533 23817 19567 23851
rect 4905 23749 4939 23783
rect 9965 23749 9999 23783
rect 23029 23749 23063 23783
rect 2513 23681 2547 23715
rect 7849 23681 7883 23715
rect 10793 23681 10827 23715
rect 1777 23613 1811 23647
rect 4813 23613 4847 23647
rect 5457 23613 5491 23647
rect 7573 23613 7607 23647
rect 9413 23613 9447 23647
rect 9689 23613 9723 23647
rect 9781 23613 9815 23647
rect 10425 23613 10459 23647
rect 10609 23613 10643 23647
rect 10701 23613 10735 23647
rect 10977 23613 11011 23647
rect 13093 23613 13127 23647
rect 13461 23613 13495 23647
rect 14105 23613 14139 23647
rect 16037 23613 16071 23647
rect 17417 23613 17451 23647
rect 18153 23613 18187 23647
rect 20085 23613 20119 23647
rect 22753 23613 22787 23647
rect 22875 23613 22909 23647
rect 23121 23613 23155 23647
rect 23949 23613 23983 23647
rect 26157 23613 26191 23647
rect 26341 23613 26375 23647
rect 26525 23613 26559 23647
rect 2780 23545 2814 23579
rect 9597 23545 9631 23579
rect 13277 23545 13311 23579
rect 13369 23545 13403 23579
rect 15301 23545 15335 23579
rect 18420 23545 18454 23579
rect 20352 23545 20386 23579
rect 24216 23545 24250 23579
rect 26433 23545 26467 23579
rect 3893 23477 3927 23511
rect 5917 23477 5951 23511
rect 11161 23477 11195 23511
rect 13645 23477 13679 23511
rect 14197 23477 14231 23511
rect 15393 23477 15427 23511
rect 16129 23477 16163 23511
rect 17509 23477 17543 23511
rect 21465 23477 21499 23511
rect 22569 23477 22603 23511
rect 25329 23477 25363 23511
rect 26709 23477 26743 23511
rect 3065 23273 3099 23307
rect 9965 23273 9999 23307
rect 10609 23273 10643 23307
rect 14933 23273 14967 23307
rect 16773 23273 16807 23307
rect 18429 23273 18463 23307
rect 23489 23273 23523 23307
rect 27445 23273 27479 23307
rect 1869 23205 1903 23239
rect 2789 23205 2823 23239
rect 18149 23205 18183 23239
rect 26332 23205 26366 23239
rect 2513 23137 2547 23171
rect 2697 23137 2731 23171
rect 2881 23137 2915 23171
rect 6653 23137 6687 23171
rect 8401 23137 8435 23171
rect 9505 23137 9539 23171
rect 10517 23137 10551 23171
rect 11428 23137 11462 23171
rect 13001 23137 13035 23171
rect 13185 23137 13219 23171
rect 13461 23137 13495 23171
rect 13737 23137 13771 23171
rect 14841 23137 14875 23171
rect 16037 23137 16071 23171
rect 16221 23137 16255 23171
rect 16589 23137 16623 23171
rect 17417 23137 17451 23171
rect 17877 23137 17911 23171
rect 18061 23137 18095 23171
rect 18245 23137 18279 23171
rect 19073 23137 19107 23171
rect 20085 23137 20119 23171
rect 20269 23137 20303 23171
rect 20361 23137 20395 23171
rect 20453 23137 20487 23171
rect 21813 23137 21847 23171
rect 23397 23137 23431 23171
rect 24225 23137 24259 23171
rect 11161 23069 11195 23103
rect 16313 23069 16347 23103
rect 16405 23069 16439 23103
rect 21557 23069 21591 23103
rect 26065 23069 26099 23103
rect 7113 23001 7147 23035
rect 13553 23001 13587 23035
rect 17233 23001 17267 23035
rect 20637 23001 20671 23035
rect 24041 23001 24075 23035
rect 1961 22933 1995 22967
rect 6837 22933 6871 22967
rect 8585 22933 8619 22967
rect 9597 22933 9631 22967
rect 12541 22933 12575 22967
rect 18889 22933 18923 22967
rect 22937 22933 22971 22967
rect 5733 22729 5767 22763
rect 10425 22729 10459 22763
rect 12173 22729 12207 22763
rect 14197 22729 14231 22763
rect 14841 22729 14875 22763
rect 26801 22729 26835 22763
rect 15669 22661 15703 22695
rect 16405 22661 16439 22695
rect 21649 22661 21683 22695
rect 24041 22593 24075 22627
rect 26065 22593 26099 22627
rect 1869 22525 1903 22559
rect 5917 22525 5951 22559
rect 6837 22525 6871 22559
rect 7021 22525 7055 22559
rect 7205 22525 7239 22559
rect 7849 22525 7883 22559
rect 8953 22525 8987 22559
rect 9873 22525 9907 22559
rect 10057 22525 10091 22559
rect 10241 22525 10275 22559
rect 11069 22525 11103 22559
rect 12081 22525 12115 22559
rect 12817 22525 12851 22559
rect 14657 22525 14691 22559
rect 15485 22525 15519 22559
rect 17325 22525 17359 22559
rect 17601 22525 17635 22559
rect 17693 22525 17727 22559
rect 18705 22525 18739 22559
rect 21097 22525 21131 22559
rect 21373 22525 21407 22559
rect 21489 22525 21523 22559
rect 22569 22525 22603 22559
rect 22937 22525 22971 22559
rect 25973 22525 26007 22559
rect 26709 22525 26743 22559
rect 2053 22457 2087 22491
rect 7113 22457 7147 22491
rect 10149 22457 10183 22491
rect 13084 22457 13118 22491
rect 16221 22457 16255 22491
rect 17509 22457 17543 22491
rect 18950 22457 18984 22491
rect 21281 22457 21315 22491
rect 22753 22457 22787 22491
rect 22845 22457 22879 22491
rect 24308 22457 24342 22491
rect 7389 22389 7423 22423
rect 7941 22389 7975 22423
rect 9045 22389 9079 22423
rect 10885 22389 10919 22423
rect 17877 22389 17911 22423
rect 20085 22389 20119 22423
rect 23121 22389 23155 22423
rect 25421 22389 25455 22423
rect 7021 22185 7055 22219
rect 11989 22185 12023 22219
rect 12449 22185 12483 22219
rect 17601 22185 17635 22219
rect 19073 22185 19107 22219
rect 25789 22185 25823 22219
rect 7665 22117 7699 22151
rect 11713 22117 11747 22151
rect 15669 22117 15703 22151
rect 21097 22117 21131 22151
rect 21281 22117 21315 22151
rect 22100 22117 22134 22151
rect 25513 22117 25547 22151
rect 26801 22117 26835 22151
rect 27537 22117 27571 22151
rect 5641 22049 5675 22083
rect 5908 22049 5942 22083
rect 7481 22049 7515 22083
rect 7757 22049 7791 22083
rect 7849 22049 7883 22083
rect 9505 22049 9539 22083
rect 9689 22049 9723 22083
rect 9777 22049 9811 22083
rect 9873 22049 9907 22083
rect 10517 22049 10551 22083
rect 11437 22049 11471 22083
rect 11621 22049 11655 22083
rect 11805 22049 11839 22083
rect 12633 22049 12667 22083
rect 13461 22049 13495 22083
rect 14749 22049 14783 22083
rect 15485 22049 15519 22083
rect 16488 22049 16522 22083
rect 18521 22049 18555 22083
rect 18705 22049 18739 22083
rect 18797 22049 18831 22083
rect 18889 22049 18923 22083
rect 19993 22049 20027 22083
rect 20177 22049 20211 22083
rect 20269 22049 20303 22083
rect 20407 22049 20441 22083
rect 21833 22049 21867 22083
rect 23673 22049 23707 22083
rect 23857 22049 23891 22083
rect 23949 22049 23983 22083
rect 24225 22049 24259 22083
rect 25237 22049 25271 22083
rect 25421 22049 25455 22083
rect 25605 22049 25639 22083
rect 26985 22049 27019 22083
rect 16221 21981 16255 22015
rect 8033 21913 8067 21947
rect 10057 21845 10091 21879
rect 10609 21845 10643 21879
rect 13553 21845 13587 21879
rect 14841 21845 14875 21879
rect 20545 21845 20579 21879
rect 23213 21845 23247 21879
rect 23673 21845 23707 21879
rect 24133 21845 24167 21879
rect 27629 21845 27663 21879
rect 2237 21641 2271 21675
rect 8217 21641 8251 21675
rect 11069 21641 11103 21675
rect 18337 21641 18371 21675
rect 23029 21641 23063 21675
rect 24225 21641 24259 21675
rect 24777 21641 24811 21675
rect 25421 21641 25455 21675
rect 9137 21573 9171 21607
rect 14086 21573 14120 21607
rect 14289 21505 14323 21539
rect 15209 21505 15243 21539
rect 19533 21505 19567 21539
rect 1685 21437 1719 21471
rect 2145 21437 2179 21471
rect 2789 21437 2823 21471
rect 4721 21437 4755 21471
rect 5365 21437 5399 21471
rect 5549 21437 5583 21471
rect 5733 21437 5767 21471
rect 6837 21437 6871 21471
rect 7104 21437 7138 21471
rect 8861 21437 8895 21471
rect 8953 21437 8987 21471
rect 9229 21437 9263 21471
rect 9689 21437 9723 21471
rect 9956 21437 9990 21471
rect 12541 21437 12575 21471
rect 13277 21437 13311 21471
rect 14151 21437 14185 21471
rect 15117 21437 15151 21471
rect 15393 21437 15427 21471
rect 15853 21437 15887 21471
rect 18061 21437 18095 21471
rect 18153 21437 18187 21471
rect 18429 21437 18463 21471
rect 18889 21437 18923 21471
rect 19800 21437 19834 21471
rect 21373 21437 21407 21471
rect 22753 21437 22787 21471
rect 22845 21437 22879 21471
rect 23121 21437 23155 21471
rect 23673 21437 23707 21471
rect 23949 21437 23983 21471
rect 24041 21437 24075 21471
rect 24685 21437 24719 21471
rect 25329 21437 25363 21471
rect 25973 21437 26007 21471
rect 26249 21437 26283 21471
rect 26341 21437 26375 21471
rect 3056 21369 3090 21403
rect 5641 21369 5675 21403
rect 13921 21369 13955 21403
rect 21465 21369 21499 21403
rect 23857 21369 23891 21403
rect 26157 21369 26191 21403
rect 1501 21301 1535 21335
rect 4169 21301 4203 21335
rect 4813 21301 4847 21335
rect 5917 21301 5951 21335
rect 8677 21301 8711 21335
rect 12725 21301 12759 21335
rect 13369 21301 13403 21335
rect 14565 21301 14599 21335
rect 17877 21301 17911 21335
rect 18981 21301 19015 21335
rect 20913 21301 20947 21335
rect 22569 21301 22603 21335
rect 26525 21301 26559 21335
rect 1961 21097 1995 21131
rect 3341 21097 3375 21131
rect 10333 21097 10367 21131
rect 11805 21097 11839 21131
rect 20177 21097 20211 21131
rect 21925 21097 21959 21131
rect 22661 21097 22695 21131
rect 25881 21097 25915 21131
rect 3065 21029 3099 21063
rect 6162 21029 6196 21063
rect 1869 20961 1903 20995
rect 2789 20961 2823 20995
rect 2973 20961 3007 20995
rect 3157 20961 3191 20995
rect 4721 20961 4755 20995
rect 4905 20961 4939 20995
rect 4997 20961 5031 20995
rect 5273 20961 5307 20995
rect 5457 20961 5491 20995
rect 8217 20961 8251 20995
rect 8309 20961 8343 20995
rect 8585 20961 8619 20995
rect 9505 20961 9539 20995
rect 10670 21029 10704 21063
rect 12449 21029 12483 21063
rect 13829 21029 13863 21063
rect 16037 21029 16071 21063
rect 17417 21029 17451 21063
rect 21741 21029 21775 21063
rect 25513 21029 25547 21063
rect 26586 21029 26620 21063
rect 12633 20961 12667 20995
rect 13093 20961 13127 20995
rect 14749 20961 14783 20995
rect 14896 20961 14930 20995
rect 17233 20961 17267 20995
rect 18153 20961 18187 20995
rect 18245 20961 18279 20995
rect 18521 20961 18555 20995
rect 20085 20961 20119 20995
rect 20729 20961 20763 20995
rect 5089 20893 5123 20927
rect 5917 20893 5951 20927
rect 10333 20893 10367 20927
rect 10425 20893 10459 20927
rect 13461 20893 13495 20927
rect 15117 20893 15151 20927
rect 13258 20825 13292 20859
rect 16221 20825 16255 20859
rect 18429 20825 18463 20859
rect 20821 20825 20855 20859
rect 21833 20961 21867 20995
rect 22569 20961 22603 20995
rect 23213 20961 23247 20995
rect 23857 20961 23891 20995
rect 25329 20961 25363 20995
rect 25605 20961 25639 20995
rect 25697 20961 25731 20995
rect 26341 20961 26375 20995
rect 7297 20757 7331 20791
rect 8033 20757 8067 20791
rect 8493 20757 8527 20791
rect 9597 20757 9631 20791
rect 13369 20757 13403 20791
rect 15025 20757 15059 20791
rect 15393 20757 15427 20791
rect 17969 20757 18003 20791
rect 21741 20757 21775 20791
rect 23305 20757 23339 20791
rect 23949 20757 23983 20791
rect 27721 20757 27755 20791
rect 3617 20553 3651 20587
rect 8585 20553 8619 20587
rect 12449 20553 12483 20587
rect 17509 20553 17543 20587
rect 19625 20553 19659 20587
rect 10701 20485 10735 20519
rect 13875 20485 13909 20519
rect 14013 20485 14047 20519
rect 16129 20485 16163 20519
rect 23857 20485 23891 20519
rect 7205 20417 7239 20451
rect 10793 20417 10827 20451
rect 14105 20417 14139 20451
rect 15761 20417 15795 20451
rect 18613 20417 18647 20451
rect 23489 20417 23523 20451
rect 1593 20349 1627 20383
rect 3525 20349 3559 20383
rect 4261 20349 4295 20383
rect 9321 20349 9355 20383
rect 10149 20349 10183 20383
rect 10241 20349 10275 20383
rect 10609 20349 10643 20383
rect 13093 20349 13127 20383
rect 13277 20349 13311 20383
rect 15301 20349 15335 20383
rect 15853 20349 15887 20383
rect 18061 20349 18095 20383
rect 18521 20349 18555 20383
rect 18889 20349 18923 20383
rect 19073 20349 19107 20383
rect 19533 20349 19567 20383
rect 20637 20349 20671 20383
rect 21005 20349 21039 20383
rect 23121 20349 23155 20383
rect 23581 20349 23615 20383
rect 23949 20349 23983 20383
rect 24133 20349 24167 20383
rect 24869 20349 24903 20383
rect 25513 20349 25547 20383
rect 25780 20349 25814 20383
rect 1860 20281 1894 20315
rect 4528 20281 4562 20315
rect 7472 20281 7506 20315
rect 12357 20281 12391 20315
rect 13737 20281 13771 20315
rect 17417 20281 17451 20315
rect 18153 20281 18187 20315
rect 20821 20281 20855 20315
rect 20913 20281 20947 20315
rect 25053 20281 25087 20315
rect 2973 20213 3007 20247
rect 5641 20213 5675 20247
rect 14381 20213 14415 20247
rect 21189 20213 21223 20247
rect 26893 20213 26927 20247
rect 2973 20009 3007 20043
rect 5825 20009 5859 20043
rect 6285 20009 6319 20043
rect 7481 20009 7515 20043
rect 8309 20009 8343 20043
rect 11989 20009 12023 20043
rect 13737 20009 13771 20043
rect 22109 20009 22143 20043
rect 2605 19941 2639 19975
rect 5549 19941 5583 19975
rect 7113 19941 7147 19975
rect 7205 19941 7239 19975
rect 18613 19941 18647 19975
rect 20996 19941 21030 19975
rect 23029 19941 23063 19975
rect 24133 19941 24167 19975
rect 1777 19873 1811 19907
rect 2421 19873 2455 19907
rect 2697 19873 2731 19907
rect 2789 19873 2823 19907
rect 5273 19873 5307 19907
rect 5457 19873 5491 19907
rect 5641 19873 5675 19907
rect 6469 19873 6503 19907
rect 6929 19873 6963 19907
rect 7297 19873 7331 19907
rect 8217 19873 8251 19907
rect 9689 19873 9723 19907
rect 9965 19873 9999 19907
rect 10425 19873 10459 19907
rect 10701 19873 10735 19907
rect 10793 19873 10827 19907
rect 11897 19873 11931 19907
rect 13093 19873 13127 19907
rect 14749 19873 14783 19907
rect 15025 19873 15059 19907
rect 16221 19873 16255 19907
rect 16488 19873 16522 19907
rect 18245 19873 18279 19907
rect 20085 19873 20119 19907
rect 22845 19873 22879 19907
rect 23121 19873 23155 19907
rect 23213 19873 23247 19907
rect 23949 19873 23983 19907
rect 26056 19873 26090 19907
rect 13461 19805 13495 19839
rect 15485 19805 15519 19839
rect 20729 19805 20763 19839
rect 25789 19805 25823 19839
rect 1961 19737 1995 19771
rect 10977 19737 11011 19771
rect 14841 19737 14875 19771
rect 20269 19737 20303 19771
rect 13231 19669 13265 19703
rect 13369 19669 13403 19703
rect 17601 19669 17635 19703
rect 23397 19669 23431 19703
rect 27169 19669 27203 19703
rect 9689 19465 9723 19499
rect 10425 19465 10459 19499
rect 14013 19465 14047 19499
rect 14381 19465 14415 19499
rect 17325 19465 17359 19499
rect 20453 19465 20487 19499
rect 13875 19397 13909 19431
rect 15025 19397 15059 19431
rect 12817 19329 12851 19363
rect 14105 19329 14139 19363
rect 17785 19329 17819 19363
rect 17877 19329 17911 19363
rect 3065 19261 3099 19295
rect 5089 19261 5123 19295
rect 5733 19261 5767 19295
rect 6837 19261 6871 19295
rect 7021 19261 7055 19295
rect 7113 19261 7147 19295
rect 7205 19261 7239 19295
rect 7389 19261 7423 19295
rect 8769 19261 8803 19295
rect 8861 19261 8895 19295
rect 9597 19261 9631 19295
rect 10241 19261 10275 19295
rect 11161 19261 11195 19295
rect 14933 19261 14967 19295
rect 15209 19261 15243 19295
rect 16129 19261 16163 19295
rect 19073 19261 19107 19295
rect 20913 19261 20947 19295
rect 21189 19261 21223 19295
rect 21281 19261 21315 19295
rect 22937 19261 22971 19295
rect 24777 19261 24811 19295
rect 26617 19261 26651 19295
rect 3332 19193 3366 19227
rect 5181 19193 5215 19227
rect 12541 19193 12575 19227
rect 13737 19193 13771 19227
rect 16221 19193 16255 19227
rect 19340 19193 19374 19227
rect 21097 19193 21131 19227
rect 23204 19193 23238 19227
rect 25022 19193 25056 19227
rect 4445 19125 4479 19159
rect 5825 19125 5859 19159
rect 7573 19125 7607 19159
rect 10977 19125 11011 19159
rect 15393 19125 15427 19159
rect 17141 19125 17175 19159
rect 17693 19125 17727 19159
rect 21465 19125 21499 19159
rect 24317 19125 24351 19159
rect 26157 19125 26191 19159
rect 4813 18921 4847 18955
rect 9689 18921 9723 18955
rect 14197 18921 14231 18955
rect 23305 18921 23339 18955
rect 26801 18921 26835 18955
rect 1501 18853 1535 18887
rect 4537 18853 4571 18887
rect 5917 18853 5951 18887
rect 2145 18785 2179 18819
rect 4261 18785 4295 18819
rect 4445 18785 4479 18819
rect 4629 18785 4663 18819
rect 5273 18785 5307 18819
rect 5365 18717 5399 18751
rect 8953 18853 8987 18887
rect 9597 18853 9631 18887
rect 13185 18853 13219 18887
rect 6009 18785 6043 18819
rect 6193 18785 6227 18819
rect 6561 18785 6595 18819
rect 7389 18785 7423 18819
rect 8033 18785 8067 18819
rect 8401 18785 8435 18819
rect 10425 18785 10459 18819
rect 11897 18785 11931 18819
rect 13001 18785 13035 18819
rect 13369 18785 13403 18819
rect 6285 18717 6319 18751
rect 6377 18717 6411 18751
rect 8309 18717 8343 18751
rect 8953 18717 8987 18751
rect 10609 18717 10643 18751
rect 7205 18649 7239 18683
rect 8493 18649 8527 18683
rect 17877 18853 17911 18887
rect 23029 18853 23063 18887
rect 25513 18853 25547 18887
rect 27537 18853 27571 18887
rect 14749 18785 14783 18819
rect 15945 18785 15979 18819
rect 16221 18785 16255 18819
rect 17141 18785 17175 18819
rect 17785 18785 17819 18819
rect 18245 18785 18279 18819
rect 18613 18785 18647 18819
rect 18797 18785 18831 18819
rect 20260 18785 20294 18819
rect 22753 18785 22787 18819
rect 22937 18785 22971 18819
rect 23121 18785 23155 18819
rect 24133 18785 24167 18819
rect 25237 18785 25271 18819
rect 25421 18785 25455 18819
rect 25605 18785 25639 18819
rect 26249 18785 26283 18819
rect 26433 18785 26467 18819
rect 26525 18785 26559 18819
rect 26617 18785 26651 18819
rect 15117 18717 15151 18751
rect 16037 18717 16071 18751
rect 16497 18717 16531 18751
rect 18337 18717 18371 18751
rect 19993 18717 20027 18751
rect 24225 18717 24259 18751
rect 15025 18649 15059 18683
rect 1593 18581 1627 18615
rect 5917 18581 5951 18615
rect 6745 18581 6779 18615
rect 8125 18581 8159 18615
rect 11989 18581 12023 18615
rect 14197 18581 14231 18615
rect 14914 18581 14948 18615
rect 15393 18581 15427 18615
rect 17233 18581 17267 18615
rect 21373 18581 21407 18615
rect 25789 18581 25823 18615
rect 27629 18581 27663 18615
rect 4537 18377 4571 18411
rect 10977 18377 11011 18411
rect 13185 18377 13219 18411
rect 19073 18377 19107 18411
rect 20545 18377 20579 18411
rect 21189 18377 21223 18411
rect 7573 18309 7607 18343
rect 14749 18309 14783 18343
rect 22661 18309 22695 18343
rect 7021 18241 7055 18275
rect 17969 18241 18003 18275
rect 25421 18241 25455 18275
rect 2145 18173 2179 18207
rect 3157 18173 3191 18207
rect 5365 18173 5399 18207
rect 5733 18173 5767 18207
rect 7389 18173 7423 18207
rect 7573 18173 7607 18207
rect 7941 18173 7975 18207
rect 9597 18173 9631 18207
rect 12081 18173 12115 18207
rect 12265 18173 12299 18207
rect 12449 18173 12483 18207
rect 13093 18173 13127 18207
rect 14657 18173 14691 18207
rect 14933 18173 14967 18207
rect 15853 18173 15887 18207
rect 17785 18173 17819 18207
rect 19993 18173 20027 18207
rect 20131 18173 20165 18207
rect 20269 18173 20303 18207
rect 20361 18173 20395 18207
rect 21005 18173 21039 18207
rect 22845 18173 22879 18207
rect 23949 18173 23983 18207
rect 1501 18105 1535 18139
rect 3424 18105 3458 18139
rect 5549 18105 5583 18139
rect 5641 18105 5675 18139
rect 9864 18105 9898 18139
rect 12357 18105 12391 18139
rect 14013 18105 14047 18139
rect 15393 18105 15427 18139
rect 18797 18105 18831 18139
rect 25666 18105 25700 18139
rect 1593 18037 1627 18071
rect 5917 18037 5951 18071
rect 12633 18037 12667 18071
rect 14105 18037 14139 18071
rect 16037 18037 16071 18071
rect 23765 18037 23799 18071
rect 26801 18037 26835 18071
rect 4813 17833 4847 17867
rect 7113 17833 7147 17867
rect 7757 17833 7791 17867
rect 8401 17833 8435 17867
rect 10517 17833 10551 17867
rect 18889 17833 18923 17867
rect 20085 17833 20119 17867
rect 4537 17765 4571 17799
rect 5978 17765 6012 17799
rect 10149 17765 10183 17799
rect 11796 17765 11830 17799
rect 15025 17765 15059 17799
rect 16313 17765 16347 17799
rect 22109 17765 22143 17799
rect 26240 17765 26274 17799
rect 1860 17697 1894 17731
rect 4307 17697 4341 17731
rect 4445 17697 4479 17731
rect 4629 17697 4663 17731
rect 7665 17697 7699 17731
rect 8309 17697 8343 17731
rect 9965 17697 9999 17731
rect 10241 17697 10275 17731
rect 10333 17697 10367 17731
rect 11529 17697 11563 17731
rect 13645 17697 13679 17731
rect 14841 17697 14875 17731
rect 15577 17697 15611 17731
rect 19073 17697 19107 17731
rect 19993 17697 20027 17731
rect 25329 17697 25363 17731
rect 25513 17697 25547 17731
rect 25973 17697 26007 17731
rect 1593 17629 1627 17663
rect 5733 17629 5767 17663
rect 13829 17561 13863 17595
rect 16497 17561 16531 17595
rect 2973 17493 3007 17527
rect 12909 17493 12943 17527
rect 15669 17493 15703 17527
rect 22201 17493 22235 17527
rect 27353 17493 27387 17527
rect 4169 17289 4203 17323
rect 4721 17289 4755 17323
rect 9137 17289 9171 17323
rect 9873 17289 9907 17323
rect 25605 17289 25639 17323
rect 5917 17221 5951 17255
rect 7113 17221 7147 17255
rect 7665 17221 7699 17255
rect 26893 17221 26927 17255
rect 1685 17153 1719 17187
rect 17877 17153 17911 17187
rect 3617 17085 3651 17119
rect 3893 17085 3927 17119
rect 3985 17085 4019 17119
rect 4629 17085 4663 17119
rect 5733 17085 5767 17119
rect 7297 17085 7331 17119
rect 7573 17085 7607 17119
rect 13553 17085 13587 17119
rect 15025 17085 15059 17119
rect 20361 17085 20395 17119
rect 20637 17085 20671 17119
rect 20729 17085 20763 17119
rect 22569 17085 22603 17119
rect 22937 17085 22971 17119
rect 25053 17085 25087 17119
rect 25329 17085 25363 17119
rect 25421 17085 25455 17119
rect 26709 17085 26743 17119
rect 1952 17017 1986 17051
rect 3801 17017 3835 17051
rect 7941 17017 7975 17051
rect 9045 17017 9079 17051
rect 9781 17017 9815 17051
rect 14381 17017 14415 17051
rect 15292 17017 15326 17051
rect 20545 17017 20579 17051
rect 22753 17017 22787 17051
rect 22845 17017 22879 17051
rect 25237 17017 25271 17051
rect 3065 16949 3099 16983
rect 13737 16949 13771 16983
rect 14473 16949 14507 16983
rect 16405 16949 16439 16983
rect 17325 16949 17359 16983
rect 17693 16949 17727 16983
rect 17785 16949 17819 16983
rect 20913 16949 20947 16983
rect 23121 16949 23155 16983
rect 1593 16745 1627 16779
rect 4353 16745 4387 16779
rect 7849 16745 7883 16779
rect 10885 16745 10919 16779
rect 11529 16745 11563 16779
rect 15301 16745 15335 16779
rect 17141 16745 17175 16779
rect 18981 16745 19015 16779
rect 21557 16745 21591 16779
rect 23949 16745 23983 16779
rect 25789 16745 25823 16779
rect 26433 16745 26467 16779
rect 2789 16677 2823 16711
rect 12633 16677 12667 16711
rect 12725 16677 12759 16711
rect 15025 16677 15059 16711
rect 16028 16677 16062 16711
rect 20444 16677 20478 16711
rect 22836 16677 22870 16711
rect 26341 16677 26375 16711
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 2697 16609 2731 16643
rect 2881 16609 2915 16643
rect 4261 16609 4295 16643
rect 6184 16609 6218 16643
rect 7757 16609 7791 16643
rect 9505 16609 9539 16643
rect 9772 16609 9806 16643
rect 11437 16609 11471 16643
rect 12449 16609 12483 16643
rect 12817 16609 12851 16643
rect 14749 16609 14783 16643
rect 14933 16609 14967 16643
rect 15117 16609 15151 16643
rect 15761 16609 15795 16643
rect 17601 16609 17635 16643
rect 17868 16609 17902 16643
rect 20177 16609 20211 16643
rect 25605 16609 25639 16643
rect 26985 16609 27019 16643
rect 5924 16541 5958 16575
rect 22569 16541 22603 16575
rect 3065 16473 3099 16507
rect 7297 16473 7331 16507
rect 13001 16405 13035 16439
rect 18981 16201 19015 16235
rect 21557 16201 21591 16235
rect 22753 16201 22787 16235
rect 25973 16201 26007 16235
rect 5917 16133 5951 16167
rect 13461 16133 13495 16167
rect 15945 16133 15979 16167
rect 17877 16133 17911 16167
rect 8493 16065 8527 16099
rect 14565 16065 14599 16099
rect 24593 16065 24627 16099
rect 2145 15997 2179 16031
rect 3617 15997 3651 16031
rect 3801 15997 3835 16031
rect 3985 15997 4019 16031
rect 4629 15997 4663 16031
rect 4997 15997 5031 16031
rect 6837 15997 6871 16031
rect 7113 15997 7147 16031
rect 7205 15997 7239 16031
rect 12081 15997 12115 16031
rect 12348 15997 12382 16031
rect 13921 15997 13955 16031
rect 3893 15929 3927 15963
rect 4813 15929 4847 15963
rect 4905 15929 4939 15963
rect 5733 15929 5767 15963
rect 7021 15929 7055 15963
rect 8738 15929 8772 15963
rect 14657 15997 14691 16031
rect 17325 15997 17359 16031
rect 17693 15997 17727 16031
rect 18889 15997 18923 16031
rect 19533 15997 19567 16031
rect 19625 15997 19659 16031
rect 23397 15997 23431 16031
rect 17509 15929 17543 15963
rect 17601 15929 17635 15963
rect 21465 15929 21499 15963
rect 22661 15929 22695 15963
rect 23581 15929 23615 15963
rect 24860 15929 24894 15963
rect 26709 15929 26743 15963
rect 4169 15861 4203 15895
rect 5181 15861 5215 15895
rect 7389 15861 7423 15895
rect 9873 15861 9907 15895
rect 14013 15861 14047 15895
rect 14565 15861 14599 15895
rect 26801 15861 26835 15895
rect 10057 15657 10091 15691
rect 23949 15657 23983 15691
rect 26617 15657 26651 15691
rect 4528 15589 4562 15623
rect 6837 15589 6871 15623
rect 7389 15589 7423 15623
rect 8585 15589 8619 15623
rect 9689 15589 9723 15623
rect 21925 15589 21959 15623
rect 27353 15589 27387 15623
rect 1409 15521 1443 15555
rect 4261 15521 4295 15555
rect 6653 15521 6687 15555
rect 8401 15521 8435 15555
rect 9505 15521 9539 15555
rect 9781 15521 9815 15555
rect 9873 15521 9907 15555
rect 10868 15521 10902 15555
rect 13369 15521 13403 15555
rect 13461 15521 13495 15555
rect 13737 15521 13771 15555
rect 15016 15521 15050 15555
rect 16865 15521 16899 15555
rect 17509 15521 17543 15555
rect 18153 15521 18187 15555
rect 18797 15521 18831 15555
rect 20260 15521 20294 15555
rect 22836 15521 22870 15555
rect 25493 15521 25527 15555
rect 27077 15521 27111 15555
rect 27261 15521 27295 15555
rect 27445 15521 27479 15555
rect 14749 15453 14783 15487
rect 19993 15453 20027 15487
rect 22569 15453 22603 15487
rect 25237 15453 25271 15487
rect 11069 15385 11103 15419
rect 16129 15385 16163 15419
rect 21373 15385 21407 15419
rect 22109 15385 22143 15419
rect 1593 15317 1627 15351
rect 5641 15317 5675 15351
rect 7481 15317 7515 15351
rect 13185 15317 13219 15351
rect 13645 15317 13679 15351
rect 16957 15317 16991 15351
rect 17601 15317 17635 15351
rect 18245 15317 18279 15351
rect 18889 15317 18923 15351
rect 27629 15317 27663 15351
rect 4353 15113 4387 15147
rect 13277 15113 13311 15147
rect 23397 15113 23431 15147
rect 24501 15113 24535 15147
rect 26893 15113 26927 15147
rect 9597 15045 9631 15079
rect 10701 15045 10735 15079
rect 15301 15045 15335 15079
rect 20269 15045 20303 15079
rect 21649 15045 21683 15079
rect 12357 14977 12391 15011
rect 14289 14977 14323 15011
rect 17785 14977 17819 15011
rect 1409 14909 1443 14943
rect 2973 14909 3007 14943
rect 3240 14909 3274 14943
rect 6837 14909 6871 14943
rect 8309 14909 8343 14943
rect 8769 14909 8803 14943
rect 9045 14909 9079 14943
rect 9321 14909 9355 14943
rect 9413 14909 9447 14943
rect 12173 14909 12207 14943
rect 13185 14909 13219 14943
rect 14749 14909 14783 14943
rect 14933 14909 14967 14943
rect 15117 14909 15151 14943
rect 17509 14909 17543 14943
rect 17601 14909 17635 14943
rect 17877 14909 17911 14943
rect 18521 14909 18555 14943
rect 19717 14909 19751 14943
rect 19901 14909 19935 14943
rect 20085 14909 20119 14943
rect 21097 14909 21131 14943
rect 21281 14909 21315 14943
rect 21465 14909 21499 14943
rect 22845 14909 22879 14943
rect 23029 14909 23063 14943
rect 23213 14909 23247 14943
rect 23949 14909 23983 14943
rect 24225 14909 24259 14943
rect 24317 14909 24351 14943
rect 25513 14909 25547 14943
rect 25780 14909 25814 14943
rect 10517 14841 10551 14875
rect 14105 14841 14139 14875
rect 15025 14841 15059 14875
rect 15853 14841 15887 14875
rect 19993 14841 20027 14875
rect 21373 14841 21407 14875
rect 23121 14841 23155 14875
rect 24133 14841 24167 14875
rect 1593 14773 1627 14807
rect 6929 14773 6963 14807
rect 15945 14773 15979 14807
rect 17325 14773 17359 14807
rect 18613 14773 18647 14807
rect 8585 14569 8619 14603
rect 22385 14569 22419 14603
rect 25881 14569 25915 14603
rect 7205 14501 7239 14535
rect 7297 14501 7331 14535
rect 9781 14501 9815 14535
rect 10517 14501 10551 14535
rect 15025 14501 15059 14535
rect 16405 14501 16439 14535
rect 21272 14501 21306 14535
rect 25605 14501 25639 14535
rect 26586 14501 26620 14535
rect 1869 14433 1903 14467
rect 4721 14433 4755 14467
rect 5917 14433 5951 14467
rect 7021 14433 7055 14467
rect 7389 14433 7423 14467
rect 8033 14433 8067 14467
rect 8217 14433 8251 14467
rect 8309 14433 8343 14467
rect 8401 14433 8435 14467
rect 9597 14433 9631 14467
rect 10241 14433 10275 14467
rect 10425 14433 10459 14467
rect 10609 14433 10643 14467
rect 11509 14433 11543 14467
rect 13645 14433 13679 14467
rect 14749 14433 14783 14467
rect 14933 14433 14967 14467
rect 15117 14433 15151 14467
rect 16221 14433 16255 14467
rect 16865 14433 16899 14467
rect 17049 14433 17083 14467
rect 17144 14433 17178 14467
rect 17233 14433 17267 14467
rect 17417 14433 17451 14467
rect 18153 14433 18187 14467
rect 20085 14433 20119 14467
rect 21005 14433 21039 14467
rect 25329 14433 25363 14467
rect 25513 14433 25547 14467
rect 25697 14433 25731 14467
rect 11253 14365 11287 14399
rect 17601 14365 17635 14399
rect 26341 14365 26375 14399
rect 2053 14297 2087 14331
rect 5181 14297 5215 14331
rect 20269 14297 20303 14331
rect 27721 14297 27755 14331
rect 4997 14229 5031 14263
rect 6009 14229 6043 14263
rect 7573 14229 7607 14263
rect 10793 14229 10827 14263
rect 12633 14229 12667 14263
rect 13737 14229 13771 14263
rect 15301 14229 15335 14263
rect 18245 14229 18279 14263
rect 8953 14025 8987 14059
rect 11161 14025 11195 14059
rect 24961 14025 24995 14059
rect 3433 13957 3467 13991
rect 13461 13957 13495 13991
rect 14289 13957 14323 13991
rect 20545 13957 20579 13991
rect 23949 13957 23983 13991
rect 26157 13957 26191 13991
rect 7573 13889 7607 13923
rect 16037 13889 16071 13923
rect 19993 13889 20027 13923
rect 1961 13821 1995 13855
rect 2145 13821 2179 13855
rect 2329 13821 2363 13855
rect 3433 13821 3467 13855
rect 3525 13821 3559 13855
rect 3709 13821 3743 13855
rect 3893 13821 3927 13855
rect 5365 13821 5399 13855
rect 5549 13821 5583 13855
rect 5733 13821 5767 13855
rect 7113 13821 7147 13855
rect 7829 13821 7863 13855
rect 9965 13821 9999 13855
rect 10609 13821 10643 13855
rect 10793 13821 10827 13855
rect 10977 13821 11011 13855
rect 12081 13821 12115 13855
rect 12337 13821 12371 13855
rect 14749 13821 14783 13855
rect 15141 13821 15175 13855
rect 17877 13821 17911 13855
rect 19809 13821 19843 13855
rect 20269 13821 20303 13855
rect 20637 13821 20671 13855
rect 20729 13821 20763 13855
rect 21373 13821 21407 13855
rect 23397 13821 23431 13855
rect 23581 13821 23615 13855
rect 23765 13821 23799 13855
rect 24409 13821 24443 13855
rect 24593 13821 24627 13855
rect 24777 13821 24811 13855
rect 25973 13821 26007 13855
rect 26617 13821 26651 13855
rect 2237 13753 2271 13787
rect 3801 13753 3835 13787
rect 5641 13753 5675 13787
rect 6929 13753 6963 13787
rect 10149 13753 10183 13787
rect 10885 13753 10919 13787
rect 14105 13753 14139 13787
rect 14933 13753 14967 13787
rect 15025 13753 15059 13787
rect 15853 13753 15887 13787
rect 18122 13753 18156 13787
rect 23673 13753 23707 13787
rect 24685 13753 24719 13787
rect 2513 13685 2547 13719
rect 4077 13685 4111 13719
rect 5917 13685 5951 13719
rect 15301 13685 15335 13719
rect 19257 13685 19291 13719
rect 21465 13685 21499 13719
rect 2881 13481 2915 13515
rect 6561 13481 6595 13515
rect 7297 13481 7331 13515
rect 8401 13481 8435 13515
rect 9689 13481 9723 13515
rect 10793 13481 10827 13515
rect 12633 13481 12667 13515
rect 16129 13481 16163 13515
rect 17693 13481 17727 13515
rect 26617 13481 26651 13515
rect 1768 13413 1802 13447
rect 5448 13413 5482 13447
rect 9597 13413 9631 13447
rect 10517 13413 10551 13447
rect 11498 13413 11532 13447
rect 15016 13413 15050 13447
rect 17325 13413 17359 13447
rect 17417 13413 17451 13447
rect 21097 13413 21131 13447
rect 22569 13413 22603 13447
rect 25482 13413 25516 13447
rect 4261 13345 4295 13379
rect 7481 13345 7515 13379
rect 7573 13345 7607 13379
rect 7849 13345 7883 13379
rect 8309 13345 8343 13379
rect 10241 13345 10275 13379
rect 10425 13345 10459 13379
rect 10609 13345 10643 13379
rect 14749 13345 14783 13379
rect 17141 13345 17175 13379
rect 17509 13345 17543 13379
rect 18245 13345 18279 13379
rect 18889 13345 18923 13379
rect 20085 13345 20119 13379
rect 21005 13345 21039 13379
rect 21465 13345 21499 13379
rect 21833 13345 21867 13379
rect 22017 13345 22051 13379
rect 22477 13345 22511 13379
rect 23213 13345 23247 13379
rect 23673 13345 23707 13379
rect 24041 13345 24075 13379
rect 24225 13345 24259 13379
rect 27077 13345 27111 13379
rect 1501 13277 1535 13311
rect 5181 13277 5215 13311
rect 11253 13277 11287 13311
rect 21557 13277 21591 13311
rect 23765 13277 23799 13311
rect 25237 13277 25271 13311
rect 7757 13209 7791 13243
rect 18981 13209 19015 13243
rect 20269 13209 20303 13243
rect 4353 13141 4387 13175
rect 18337 13141 18371 13175
rect 23305 13141 23339 13175
rect 4261 12937 4295 12971
rect 8217 12937 8251 12971
rect 8769 12937 8803 12971
rect 15945 12937 15979 12971
rect 10977 12869 11011 12903
rect 17785 12869 17819 12903
rect 2881 12801 2915 12835
rect 6837 12801 6871 12835
rect 12173 12801 12207 12835
rect 23029 12801 23063 12835
rect 1409 12733 1443 12767
rect 2053 12733 2087 12767
rect 3148 12733 3182 12767
rect 4721 12733 4755 12767
rect 5365 12733 5399 12767
rect 5549 12733 5583 12767
rect 5641 12733 5675 12767
rect 5733 12733 5767 12767
rect 8677 12733 8711 12767
rect 9505 12733 9539 12767
rect 9689 12733 9723 12767
rect 9781 12733 9815 12767
rect 9873 12733 9907 12767
rect 10057 12733 10091 12767
rect 12081 12733 12115 12767
rect 13829 12733 13863 12767
rect 14565 12733 14599 12767
rect 14832 12733 14866 12767
rect 17325 12733 17359 12767
rect 17509 12733 17543 12767
rect 17601 12733 17635 12767
rect 17877 12733 17911 12767
rect 18337 12733 18371 12767
rect 19625 12733 19659 12767
rect 20269 12733 20303 12767
rect 25145 12733 25179 12767
rect 7082 12665 7116 12699
rect 10793 12665 10827 12699
rect 19809 12665 19843 12699
rect 20536 12665 20570 12699
rect 23296 12665 23330 12699
rect 25412 12665 25446 12699
rect 2237 12597 2271 12631
rect 4813 12597 4847 12631
rect 5917 12597 5951 12631
rect 10241 12597 10275 12631
rect 14013 12597 14047 12631
rect 17325 12597 17359 12631
rect 18521 12597 18555 12631
rect 21649 12597 21683 12631
rect 24409 12597 24443 12631
rect 26525 12597 26559 12631
rect 11713 12393 11747 12427
rect 14933 12393 14967 12427
rect 17233 12393 17267 12427
rect 18429 12393 18463 12427
rect 22017 12393 22051 12427
rect 22569 12393 22603 12427
rect 23673 12393 23707 12427
rect 24225 12393 24259 12427
rect 25789 12393 25823 12427
rect 7205 12325 7239 12359
rect 10057 12325 10091 12359
rect 10977 12325 11011 12359
rect 23305 12325 23339 12359
rect 23397 12325 23431 12359
rect 25421 12325 25455 12359
rect 26801 12325 26835 12359
rect 27537 12325 27571 12359
rect 1961 12257 1995 12291
rect 2228 12257 2262 12291
rect 4537 12257 4571 12291
rect 4721 12257 4755 12291
rect 4905 12257 4939 12291
rect 5089 12257 5123 12291
rect 6101 12257 6135 12291
rect 6285 12257 6319 12291
rect 6561 12257 6595 12291
rect 9781 12257 9815 12291
rect 9965 12257 9999 12291
rect 10149 12257 10183 12291
rect 11621 12257 11655 12291
rect 12449 12257 12483 12291
rect 13001 12257 13035 12291
rect 14841 12257 14875 12291
rect 15669 12257 15703 12291
rect 15761 12257 15795 12291
rect 16037 12257 16071 12291
rect 16497 12257 16531 12291
rect 16681 12257 16715 12291
rect 16865 12257 16899 12291
rect 17049 12257 17083 12291
rect 17693 12257 17727 12291
rect 18337 12257 18371 12291
rect 20904 12257 20938 12291
rect 22477 12257 22511 12291
rect 23121 12257 23155 12291
rect 23489 12257 23523 12291
rect 24133 12257 24167 12291
rect 25237 12257 25271 12291
rect 25513 12257 25547 12291
rect 25605 12257 25639 12291
rect 27721 12257 27755 12291
rect 4813 12189 4847 12223
rect 15485 12189 15519 12223
rect 16773 12189 16807 12223
rect 20637 12189 20671 12223
rect 5273 12121 5307 12155
rect 5825 12121 5859 12155
rect 6377 12121 6411 12155
rect 17785 12121 17819 12155
rect 3341 12053 3375 12087
rect 7297 12053 7331 12087
rect 10333 12053 10367 12087
rect 11069 12053 11103 12087
rect 12265 12053 12299 12087
rect 13093 12053 13127 12087
rect 15945 12053 15979 12087
rect 26893 12053 26927 12087
rect 21189 11849 21223 11883
rect 24869 11849 24903 11883
rect 25421 11849 25455 11883
rect 3709 11781 3743 11815
rect 4261 11781 4295 11815
rect 5549 11781 5583 11815
rect 8677 11781 8711 11815
rect 10701 11781 10735 11815
rect 13829 11781 13863 11815
rect 13369 11713 13403 11747
rect 13921 11713 13955 11747
rect 1501 11645 1535 11679
rect 2145 11645 2179 11679
rect 3157 11645 3191 11679
rect 3433 11645 3467 11679
rect 3525 11645 3559 11679
rect 4169 11645 4203 11679
rect 5733 11645 5767 11679
rect 6929 11645 6963 11679
rect 9321 11645 9355 11679
rect 9588 11645 9622 11679
rect 13185 11645 13219 11679
rect 13645 11645 13679 11679
rect 14013 11645 14047 11679
rect 15761 11645 15795 11679
rect 15945 11645 15979 11679
rect 17325 11645 17359 11679
rect 19441 11645 19475 11679
rect 20085 11645 20119 11679
rect 20637 11645 20671 11679
rect 21005 11645 21039 11679
rect 23213 11645 23247 11679
rect 24041 11645 24075 11679
rect 24777 11645 24811 11679
rect 25605 11645 25639 11679
rect 26065 11645 26099 11679
rect 26433 11645 26467 11679
rect 1685 11577 1719 11611
rect 3341 11577 3375 11611
rect 8493 11577 8527 11611
rect 12173 11577 12207 11611
rect 12357 11577 12391 11611
rect 16129 11577 16163 11611
rect 17570 11577 17604 11611
rect 20821 11577 20855 11611
rect 20913 11577 20947 11611
rect 26249 11577 26283 11611
rect 26341 11577 26375 11611
rect 7021 11509 7055 11543
rect 18705 11509 18739 11543
rect 19257 11509 19291 11543
rect 19901 11509 19935 11543
rect 23305 11509 23339 11543
rect 23857 11509 23891 11543
rect 26617 11509 26651 11543
rect 6929 11305 6963 11339
rect 13737 11305 13771 11339
rect 17325 11305 17359 11339
rect 18245 11305 18279 11339
rect 21097 11305 21131 11339
rect 27721 11305 27755 11339
rect 4537 11237 4571 11271
rect 12173 11237 12207 11271
rect 14933 11237 14967 11271
rect 16957 11237 16991 11271
rect 17049 11237 17083 11271
rect 20821 11237 20855 11271
rect 22477 11237 22511 11271
rect 22569 11237 22603 11271
rect 23397 11237 23431 11271
rect 25605 11237 25639 11271
rect 26608 11237 26642 11271
rect 4261 11169 4295 11203
rect 4445 11169 4479 11203
rect 4629 11169 4663 11203
rect 5733 11169 5767 11203
rect 7113 11169 7147 11203
rect 8125 11169 8159 11203
rect 8493 11169 8527 11203
rect 10324 11169 10358 11203
rect 11897 11169 11931 11203
rect 12081 11169 12115 11203
rect 12265 11169 12299 11203
rect 12909 11169 12943 11203
rect 13637 11169 13671 11203
rect 14749 11169 14783 11203
rect 15025 11169 15059 11203
rect 15117 11169 15151 11203
rect 15761 11169 15795 11203
rect 16773 11169 16807 11203
rect 17141 11169 17175 11203
rect 18061 11169 18095 11203
rect 18889 11169 18923 11203
rect 20545 11169 20579 11203
rect 20729 11169 20763 11203
rect 20913 11169 20947 11203
rect 22293 11169 22327 11203
rect 22661 11169 22695 11203
rect 23305 11169 23339 11203
rect 23765 11169 23799 11203
rect 24133 11169 24167 11203
rect 24317 11169 24351 11203
rect 25329 11169 25363 11203
rect 25513 11169 25547 11203
rect 25697 11169 25731 11203
rect 26341 11169 26375 11203
rect 8401 11101 8435 11135
rect 10057 11101 10091 11135
rect 23857 11101 23891 11135
rect 5825 11033 5859 11067
rect 13093 11033 13127 11067
rect 15945 11033 15979 11067
rect 4813 10965 4847 10999
rect 8217 10965 8251 10999
rect 8585 10965 8619 10999
rect 11437 10965 11471 10999
rect 12449 10965 12483 10999
rect 15301 10965 15335 10999
rect 18981 10965 19015 10999
rect 22845 10965 22879 10999
rect 25881 10965 25915 10999
rect 10149 10761 10183 10795
rect 11161 10761 11195 10795
rect 13461 10761 13495 10795
rect 24961 10761 24995 10795
rect 8309 10693 8343 10727
rect 2697 10625 2731 10659
rect 4997 10625 5031 10659
rect 5089 10625 5123 10659
rect 7021 10625 7055 10659
rect 8769 10625 8803 10659
rect 12081 10625 12115 10659
rect 14657 10625 14691 10659
rect 18153 10625 18187 10659
rect 18245 10625 18279 10659
rect 19625 10625 19659 10659
rect 1869 10557 1903 10591
rect 4721 10557 4755 10591
rect 4905 10557 4939 10591
rect 5273 10557 5307 10591
rect 7297 10557 7331 10591
rect 7573 10557 7607 10591
rect 7941 10557 7975 10591
rect 10609 10557 10643 10591
rect 10793 10557 10827 10591
rect 10977 10557 11011 10591
rect 14924 10557 14958 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 18429 10557 18463 10591
rect 22753 10557 22787 10591
rect 24869 10557 24903 10591
rect 25513 10557 25547 10591
rect 25780 10557 25814 10591
rect 2964 10489 2998 10523
rect 5457 10489 5491 10523
rect 9036 10489 9070 10523
rect 10885 10489 10919 10523
rect 12348 10489 12382 10523
rect 14013 10489 14047 10523
rect 19892 10489 19926 10523
rect 23020 10489 23054 10523
rect 1961 10421 1995 10455
rect 4077 10421 4111 10455
rect 14105 10421 14139 10455
rect 16037 10421 16071 10455
rect 18613 10421 18647 10455
rect 21005 10421 21039 10455
rect 24133 10421 24167 10455
rect 26893 10421 26927 10455
rect 2881 10217 2915 10251
rect 5641 10217 5675 10251
rect 10057 10217 10091 10251
rect 17601 10217 17635 10251
rect 18153 10217 18187 10251
rect 21373 10217 21407 10251
rect 23673 10217 23707 10251
rect 24225 10217 24259 10251
rect 26709 10217 26743 10251
rect 4528 10149 4562 10183
rect 10609 10149 10643 10183
rect 12081 10149 12115 10183
rect 22560 10149 22594 10183
rect 27537 10149 27571 10183
rect 27721 10149 27755 10183
rect 1768 10081 1802 10115
rect 4261 10081 4295 10115
rect 6357 10081 6391 10115
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 9781 10081 9815 10115
rect 9919 10081 9953 10115
rect 10517 10081 10551 10115
rect 11897 10081 11931 10115
rect 12173 10081 12207 10115
rect 12265 10081 12299 10115
rect 16221 10081 16255 10115
rect 16488 10081 16522 10115
rect 18337 10081 18371 10115
rect 18429 10081 18463 10115
rect 18705 10081 18739 10115
rect 19993 10081 20027 10115
rect 20260 10081 20294 10115
rect 22293 10081 22327 10115
rect 24133 10081 24167 10115
rect 25329 10081 25363 10115
rect 25596 10081 25630 10115
rect 1501 10013 1535 10047
rect 6101 10013 6135 10047
rect 7481 9877 7515 9911
rect 12449 9877 12483 9911
rect 18613 9877 18647 9911
rect 5917 9673 5951 9707
rect 10057 9605 10091 9639
rect 13829 9605 13863 9639
rect 17325 9605 17359 9639
rect 19257 9605 19291 9639
rect 20729 9605 20763 9639
rect 2053 9537 2087 9571
rect 6837 9537 6871 9571
rect 12449 9537 12483 9571
rect 17877 9537 17911 9571
rect 21281 9537 21315 9571
rect 23029 9537 23063 9571
rect 23305 9537 23339 9571
rect 1409 9469 1443 9503
rect 3985 9469 4019 9503
rect 4261 9469 4295 9503
rect 4353 9469 4387 9503
rect 5365 9469 5399 9503
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 8677 9469 8711 9503
rect 9321 9469 9355 9503
rect 10241 9469 10275 9503
rect 10977 9469 11011 9503
rect 12705 9469 12739 9503
rect 14473 9469 14507 9503
rect 18705 9469 18739 9503
rect 18981 9469 19015 9503
rect 19165 9469 19199 9503
rect 19533 9469 19567 9503
rect 19717 9469 19751 9503
rect 20177 9469 20211 9503
rect 20545 9469 20579 9503
rect 21189 9469 21223 9503
rect 22937 9469 22971 9503
rect 23397 9469 23431 9503
rect 23765 9469 23799 9503
rect 23949 9469 23983 9503
rect 24869 9469 24903 9503
rect 26709 9469 26743 9503
rect 2320 9401 2354 9435
rect 4169 9401 4203 9435
rect 5549 9401 5583 9435
rect 7082 9401 7116 9435
rect 14657 9401 14691 9435
rect 17785 9401 17819 9435
rect 20361 9401 20395 9435
rect 20453 9401 20487 9435
rect 25136 9401 25170 9435
rect 1593 9333 1627 9367
rect 3433 9333 3467 9367
rect 4537 9333 4571 9367
rect 8217 9333 8251 9367
rect 8769 9333 8803 9367
rect 9413 9333 9447 9367
rect 11069 9333 11103 9367
rect 17693 9333 17727 9367
rect 26249 9333 26283 9367
rect 2697 9129 2731 9163
rect 4445 9129 4479 9163
rect 5181 9129 5215 9163
rect 6929 9129 6963 9163
rect 16773 9129 16807 9163
rect 20545 9129 20579 9163
rect 23305 9129 23339 9163
rect 24225 9129 24259 9163
rect 25789 9129 25823 9163
rect 26985 9129 27019 9163
rect 2421 9061 2455 9095
rect 6653 9061 6687 9095
rect 9689 9061 9723 9095
rect 10977 9061 11011 9095
rect 12725 9061 12759 9095
rect 15025 9061 15059 9095
rect 17693 9061 17727 9095
rect 20177 9061 20211 9095
rect 20269 9061 20303 9095
rect 22937 9061 22971 9095
rect 25421 9061 25455 9095
rect 25513 9061 25547 9095
rect 1409 8993 1443 9027
rect 2145 8993 2179 9027
rect 2329 8993 2363 9027
rect 2513 8993 2547 9027
rect 3157 8993 3191 9027
rect 4353 8993 4387 9027
rect 5089 8993 5123 9027
rect 5917 8993 5951 9027
rect 6377 8993 6411 9027
rect 6561 8993 6595 9027
rect 6745 8993 6779 9027
rect 7573 8993 7607 9027
rect 8033 8993 8067 9027
rect 8401 8993 8435 9027
rect 9505 8993 9539 9027
rect 9789 8993 9823 9027
rect 9919 8993 9953 9027
rect 10885 8993 10919 9027
rect 11069 8993 11103 9027
rect 11345 8993 11379 9027
rect 11713 8993 11747 9027
rect 11897 8993 11931 9027
rect 13369 8993 13403 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15117 8993 15151 9027
rect 16589 8993 16623 9027
rect 18429 8993 18463 9027
rect 19993 8993 20027 9027
rect 20361 8993 20395 9027
rect 22753 8993 22787 9027
rect 23029 8993 23063 9027
rect 23121 8993 23155 9027
rect 24133 8993 24167 9027
rect 25237 8993 25271 9027
rect 25629 8993 25663 9027
rect 26801 8993 26835 9027
rect 27537 8993 27571 9027
rect 3249 8925 3283 8959
rect 7757 8925 7791 8959
rect 8309 8925 8343 8959
rect 5733 8857 5767 8891
rect 8217 8857 8251 8891
rect 17877 8857 17911 8891
rect 27721 8857 27755 8891
rect 10057 8789 10091 8823
rect 12817 8789 12851 8823
rect 13553 8789 13587 8823
rect 15301 8789 15335 8823
rect 18521 8789 18555 8823
rect 2881 8585 2915 8619
rect 4077 8585 4111 8619
rect 4353 8585 4387 8619
rect 7665 8585 7699 8619
rect 9597 8585 9631 8619
rect 15761 8585 15795 8619
rect 18245 8585 18279 8619
rect 20177 8585 20211 8619
rect 25145 8585 25179 8619
rect 10793 8517 10827 8551
rect 13921 8517 13955 8551
rect 17601 8517 17635 8551
rect 26157 8517 26191 8551
rect 10241 8449 10275 8483
rect 2329 8381 2363 8415
rect 2513 8381 2547 8415
rect 2697 8381 2731 8415
rect 3893 8381 3927 8415
rect 6837 8381 6871 8415
rect 7573 8381 7607 8415
rect 8217 8381 8251 8415
rect 8484 8381 8518 8415
rect 10057 8381 10091 8415
rect 10517 8381 10551 8415
rect 10885 8381 10919 8415
rect 10977 8381 11011 8415
rect 12081 8381 12115 8415
rect 12357 8381 12391 8415
rect 12449 8381 12483 8415
rect 13369 8381 13403 8415
rect 13645 8381 13679 8415
rect 13737 8381 13771 8415
rect 14381 8381 14415 8415
rect 14637 8381 14671 8415
rect 17417 8381 17451 8415
rect 18153 8381 18187 8415
rect 18797 8381 18831 8415
rect 19064 8381 19098 8415
rect 20729 8381 20763 8415
rect 21557 8381 21591 8415
rect 22753 8381 22787 8415
rect 24133 8381 24167 8415
rect 24593 8381 24627 8415
rect 24869 8381 24903 8415
rect 24961 8381 24995 8415
rect 25605 8381 25639 8415
rect 25881 8381 25915 8415
rect 25973 8381 26007 8415
rect 26709 8381 26743 8415
rect 2605 8313 2639 8347
rect 12265 8313 12299 8347
rect 13553 8313 13587 8347
rect 24777 8313 24811 8347
rect 25789 8313 25823 8347
rect 6929 8245 6963 8279
rect 12633 8245 12667 8279
rect 20821 8245 20855 8279
rect 21373 8245 21407 8279
rect 22845 8245 22879 8279
rect 23949 8245 23983 8279
rect 26893 8245 26927 8279
rect 1593 8041 1627 8075
rect 7849 8041 7883 8075
rect 9873 8041 9907 8075
rect 13737 8041 13771 8075
rect 17049 8041 17083 8075
rect 20361 8041 20395 8075
rect 21189 8041 21223 8075
rect 23397 8041 23431 8075
rect 27353 8041 27387 8075
rect 4721 7973 4755 8007
rect 5724 7973 5758 8007
rect 12624 7973 12658 8007
rect 15016 7973 15050 8007
rect 1409 7905 1443 7939
rect 2145 7905 2179 7939
rect 4445 7905 4479 7939
rect 4629 7905 4663 7939
rect 4813 7905 4847 7939
rect 5457 7905 5491 7939
rect 7297 7905 7331 7939
rect 7481 7905 7515 7939
rect 7573 7905 7607 7939
rect 7665 7905 7699 7939
rect 10057 7905 10091 7939
rect 10517 7905 10551 7939
rect 10784 7905 10818 7939
rect 12357 7905 12391 7939
rect 14749 7905 14783 7939
rect 16589 7905 16623 7939
rect 17509 7905 17543 7939
rect 17693 7905 17727 7939
rect 17785 7905 17819 7939
rect 17877 7905 17911 7939
rect 18521 7905 18555 7939
rect 18705 7905 18739 7939
rect 18797 7905 18831 7939
rect 18889 7905 18923 7939
rect 21741 7973 21775 8007
rect 26240 7973 26274 8007
rect 20453 7905 20487 7939
rect 20637 7905 20671 7939
rect 20867 7905 20901 7939
rect 21005 7905 21039 7939
rect 21649 7905 21683 7939
rect 22661 7905 22695 7939
rect 22845 7905 22879 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 24133 7905 24167 7939
rect 25237 7905 25271 7939
rect 20361 7837 20395 7871
rect 20729 7837 20763 7871
rect 22937 7837 22971 7871
rect 24225 7837 24259 7871
rect 25973 7837 26007 7871
rect 6837 7769 6871 7803
rect 4997 7701 5031 7735
rect 11897 7701 11931 7735
rect 16129 7701 16163 7735
rect 16865 7701 16899 7735
rect 18061 7701 18095 7735
rect 19073 7701 19107 7735
rect 20361 7701 20395 7735
rect 25329 7701 25363 7735
rect 1593 7497 1627 7531
rect 3801 7497 3835 7531
rect 5825 7497 5859 7531
rect 10609 7497 10643 7531
rect 12173 7497 12207 7531
rect 16313 7497 16347 7531
rect 19717 7497 19751 7531
rect 20085 7497 20119 7531
rect 23305 7497 23339 7531
rect 26249 7497 26283 7531
rect 3985 7429 4019 7463
rect 7297 7429 7331 7463
rect 11069 7429 11103 7463
rect 4445 7361 4479 7395
rect 6837 7361 6871 7395
rect 17693 7361 17727 7395
rect 22845 7361 22879 7395
rect 22937 7361 22971 7395
rect 1501 7293 1535 7327
rect 2145 7293 2179 7327
rect 2329 7293 2363 7327
rect 2513 7293 2547 7327
rect 3547 7293 3581 7327
rect 4712 7293 4746 7327
rect 7021 7293 7055 7327
rect 7113 7293 7147 7327
rect 7389 7293 7423 7327
rect 7849 7293 7883 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 11161 7293 11195 7327
rect 12081 7293 12115 7327
rect 12725 7293 12759 7327
rect 16221 7293 16255 7327
rect 17960 7293 17994 7327
rect 19625 7293 19659 7327
rect 21097 7293 21131 7327
rect 21281 7293 21315 7327
rect 21465 7293 21499 7327
rect 22569 7293 22603 7327
rect 22753 7293 22787 7327
rect 23121 7293 23155 7327
rect 23857 7293 23891 7327
rect 24133 7293 24167 7327
rect 24225 7293 24259 7327
rect 24869 7293 24903 7327
rect 2421 7225 2455 7259
rect 12817 7225 12851 7259
rect 21373 7225 21407 7259
rect 24041 7225 24075 7259
rect 25114 7225 25148 7259
rect 2697 7157 2731 7191
rect 7941 7157 7975 7191
rect 19073 7157 19107 7191
rect 21649 7157 21683 7191
rect 24409 7157 24443 7191
rect 11437 6953 11471 6987
rect 2044 6885 2078 6919
rect 4537 6885 4571 6919
rect 5733 6885 5767 6919
rect 11161 6885 11195 6919
rect 20269 6885 20303 6919
rect 22906 6885 22940 6919
rect 25513 6885 25547 6919
rect 4261 6817 4295 6851
rect 4445 6817 4479 6851
rect 4629 6817 4663 6851
rect 5549 6817 5583 6851
rect 6193 6817 6227 6851
rect 7389 6817 7423 6851
rect 7481 6817 7515 6851
rect 7757 6817 7791 6851
rect 10885 6817 10919 6851
rect 11069 6817 11103 6851
rect 11253 6817 11287 6851
rect 12173 6817 12207 6851
rect 15761 6817 15795 6851
rect 16028 6817 16062 6851
rect 18061 6817 18095 6851
rect 18705 6817 18739 6851
rect 20177 6817 20211 6851
rect 20821 6817 20855 6851
rect 21088 6817 21122 6851
rect 25237 6817 25271 6851
rect 25421 6817 25455 6851
rect 25605 6817 25639 6851
rect 26505 6817 26539 6851
rect 1777 6749 1811 6783
rect 7205 6749 7239 6783
rect 18153 6749 18187 6783
rect 22661 6749 22695 6783
rect 26249 6749 26283 6783
rect 7665 6681 7699 6715
rect 18797 6681 18831 6715
rect 25789 6681 25823 6715
rect 27629 6681 27663 6715
rect 3157 6613 3191 6647
rect 4813 6613 4847 6647
rect 6285 6613 6319 6647
rect 12265 6613 12299 6647
rect 17141 6613 17175 6647
rect 22201 6613 22235 6647
rect 24041 6613 24075 6647
rect 1593 6409 1627 6443
rect 4261 6409 4295 6443
rect 5641 6409 5675 6443
rect 8401 6409 8435 6443
rect 9413 6409 9447 6443
rect 13093 6409 13127 6443
rect 16405 6409 16439 6443
rect 17693 6409 17727 6443
rect 21097 6409 21131 6443
rect 23857 6409 23891 6443
rect 24409 6409 24443 6443
rect 26801 6409 26835 6443
rect 4997 6273 5031 6307
rect 12725 6273 12759 6307
rect 19349 6273 19383 6307
rect 23397 6273 23431 6307
rect 1409 6205 1443 6239
rect 2881 6205 2915 6239
rect 3148 6205 3182 6239
rect 4813 6205 4847 6239
rect 5457 6205 5491 6239
rect 8108 6205 8142 6239
rect 8217 6205 8251 6239
rect 8493 6205 8527 6239
rect 8953 6205 8987 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 9505 6205 9539 6239
rect 12633 6205 12667 6239
rect 12817 6205 12851 6239
rect 12909 6205 12943 6239
rect 13185 6205 13219 6239
rect 14013 6205 14047 6239
rect 14197 6205 14231 6239
rect 14381 6205 14415 6239
rect 15393 6205 15427 6239
rect 15853 6205 15887 6239
rect 16221 6205 16255 6239
rect 17509 6205 17543 6239
rect 18337 6205 18371 6239
rect 20545 6205 20579 6239
rect 20821 6205 20855 6239
rect 20913 6205 20947 6239
rect 23121 6205 23155 6239
rect 23305 6205 23339 6239
rect 23489 6205 23523 6239
rect 23673 6205 23707 6239
rect 24317 6205 24351 6239
rect 26709 6205 26743 6239
rect 14289 6137 14323 6171
rect 16037 6137 16071 6171
rect 16129 6137 16163 6171
rect 19165 6137 19199 6171
rect 20729 6137 20763 6171
rect 7941 6069 7975 6103
rect 8953 6069 8987 6103
rect 14565 6069 14599 6103
rect 15209 6069 15243 6103
rect 18429 6069 18463 6103
rect 24777 6069 24811 6103
rect 4353 5865 4387 5899
rect 8585 5865 8619 5899
rect 10057 5865 10091 5899
rect 10609 5865 10643 5899
rect 12817 5865 12851 5899
rect 14841 5865 14875 5899
rect 16865 5865 16899 5899
rect 21557 5865 21591 5899
rect 23029 5865 23063 5899
rect 7472 5797 7506 5831
rect 9781 5797 9815 5831
rect 18889 5797 18923 5831
rect 19073 5797 19107 5831
rect 23765 5797 23799 5831
rect 27537 5797 27571 5831
rect 27721 5797 27755 5831
rect 4261 5729 4295 5763
rect 7205 5729 7239 5763
rect 9505 5729 9539 5763
rect 9689 5729 9723 5763
rect 9873 5729 9907 5763
rect 10517 5729 10551 5763
rect 11253 5729 11287 5763
rect 11437 5729 11471 5763
rect 11529 5729 11563 5763
rect 11667 5729 11701 5763
rect 13001 5729 13035 5763
rect 13093 5729 13127 5763
rect 13369 5729 13403 5763
rect 14749 5729 14783 5763
rect 15752 5729 15786 5763
rect 17509 5729 17543 5763
rect 20177 5729 20211 5763
rect 21097 5729 21131 5763
rect 22569 5729 22603 5763
rect 23489 5729 23523 5763
rect 23673 5729 23707 5763
rect 23857 5729 23891 5763
rect 13277 5661 13311 5695
rect 15485 5661 15519 5695
rect 17785 5661 17819 5695
rect 11805 5525 11839 5559
rect 19993 5525 20027 5559
rect 21189 5525 21223 5559
rect 22845 5525 22879 5559
rect 24041 5525 24075 5559
rect 3525 5321 3559 5355
rect 7205 5321 7239 5355
rect 25145 5321 25179 5355
rect 7849 5253 7883 5287
rect 10793 5253 10827 5287
rect 15117 5253 15151 5287
rect 16405 5253 16439 5287
rect 21557 5253 21591 5287
rect 2145 5185 2179 5219
rect 8401 5185 8435 5219
rect 17601 5185 17635 5219
rect 19073 5185 19107 5219
rect 23765 5185 23799 5219
rect 1409 5117 1443 5151
rect 7113 5117 7147 5151
rect 7757 5117 7791 5151
rect 10241 5117 10275 5151
rect 10425 5117 10459 5151
rect 10609 5117 10643 5151
rect 12081 5117 12115 5151
rect 12449 5117 12483 5151
rect 13093 5117 13127 5151
rect 15025 5117 15059 5151
rect 15853 5117 15887 5151
rect 16221 5117 16255 5151
rect 17417 5117 17451 5151
rect 18061 5117 18095 5151
rect 18429 5117 18463 5151
rect 21465 5117 21499 5151
rect 22661 5117 22695 5151
rect 22937 5117 22971 5151
rect 23029 5117 23063 5151
rect 26709 5117 26743 5151
rect 2412 5049 2446 5083
rect 8668 5049 8702 5083
rect 10517 5049 10551 5083
rect 12265 5049 12299 5083
rect 12357 5049 12391 5083
rect 13360 5049 13394 5083
rect 16037 5049 16071 5083
rect 16129 5049 16163 5083
rect 18245 5049 18279 5083
rect 18337 5049 18371 5083
rect 19340 5049 19374 5083
rect 22845 5049 22879 5083
rect 24032 5049 24066 5083
rect 1593 4981 1627 5015
rect 9781 4981 9815 5015
rect 12633 4981 12667 5015
rect 14473 4981 14507 5015
rect 18613 4981 18647 5015
rect 20453 4981 20487 5015
rect 23213 4981 23247 5015
rect 26893 4981 26927 5015
rect 6837 4777 6871 4811
rect 8493 4777 8527 4811
rect 10149 4777 10183 4811
rect 12449 4777 12483 4811
rect 13461 4777 13495 4811
rect 20545 4777 20579 4811
rect 21005 4777 21039 4811
rect 24225 4777 24259 4811
rect 1685 4709 1719 4743
rect 2605 4709 2639 4743
rect 9781 4709 9815 4743
rect 11336 4709 11370 4743
rect 13093 4709 13127 4743
rect 15016 4709 15050 4743
rect 17049 4709 17083 4743
rect 17960 4709 17994 4743
rect 20269 4709 20303 4743
rect 23112 4709 23146 4743
rect 27537 4709 27571 4743
rect 2329 4641 2363 4675
rect 2513 4641 2547 4675
rect 2697 4641 2731 4675
rect 5069 4641 5103 4675
rect 6745 4641 6779 4675
rect 8401 4641 8435 4675
rect 9597 4641 9631 4675
rect 9873 4641 9907 4675
rect 9965 4641 9999 4675
rect 11069 4641 11103 4675
rect 12909 4641 12943 4675
rect 13185 4641 13219 4675
rect 13277 4641 13311 4675
rect 14749 4641 14783 4675
rect 17693 4641 17727 4675
rect 19993 4641 20027 4675
rect 20177 4641 20211 4675
rect 20361 4641 20395 4675
rect 21189 4641 21223 4675
rect 21833 4641 21867 4675
rect 25421 4641 25455 4675
rect 26157 4641 26191 4675
rect 26801 4641 26835 4675
rect 4813 4573 4847 4607
rect 22845 4573 22879 4607
rect 27721 4573 27755 4607
rect 2881 4505 2915 4539
rect 17233 4505 17267 4539
rect 21649 4505 21683 4539
rect 26985 4505 27019 4539
rect 1777 4437 1811 4471
rect 6193 4437 6227 4471
rect 16129 4437 16163 4471
rect 19073 4437 19107 4471
rect 25237 4437 25271 4471
rect 26341 4437 26375 4471
rect 2513 4233 2547 4267
rect 4905 4233 4939 4267
rect 10333 4233 10367 4267
rect 13461 4233 13495 4267
rect 14657 4233 14691 4267
rect 20361 4165 20395 4199
rect 8953 4097 8987 4131
rect 11069 4097 11103 4131
rect 12081 4097 12115 4131
rect 14013 4097 14047 4131
rect 22661 4097 22695 4131
rect 23305 4097 23339 4131
rect 2697 4029 2731 4063
rect 3157 4029 3191 4063
rect 4353 4029 4387 4063
rect 4629 4029 4663 4063
rect 4721 4029 4755 4063
rect 5365 4029 5399 4063
rect 5733 4029 5767 4063
rect 9220 4029 9254 4063
rect 12348 4029 12382 4063
rect 13921 4029 13955 4063
rect 14565 4029 14599 4063
rect 15209 4029 15243 4063
rect 17325 4029 17359 4063
rect 17969 4029 18003 4063
rect 18337 4029 18371 4063
rect 18981 4029 19015 4063
rect 19237 4029 19271 4063
rect 21189 4029 21223 4063
rect 22569 4029 22603 4063
rect 23213 4029 23247 4063
rect 24041 4029 24075 4063
rect 24869 4029 24903 4063
rect 25973 4029 26007 4063
rect 1869 3961 1903 3995
rect 4537 3961 4571 3995
rect 5549 3961 5583 3995
rect 5641 3961 5675 3995
rect 10885 3961 10919 3995
rect 16221 3961 16255 3995
rect 17417 3961 17451 3995
rect 18153 3961 18187 3995
rect 18245 3961 18279 3995
rect 26709 3961 26743 3995
rect 26893 3961 26927 3995
rect 1961 3893 1995 3927
rect 3341 3893 3375 3927
rect 5917 3893 5951 3927
rect 16313 3893 16347 3927
rect 18521 3893 18555 3927
rect 23857 3893 23891 3927
rect 25053 3893 25087 3927
rect 26157 3893 26191 3927
rect 6929 3689 6963 3723
rect 18981 3689 19015 3723
rect 5816 3621 5850 3655
rect 10241 3621 10275 3655
rect 13093 3621 13127 3655
rect 14933 3621 14967 3655
rect 20913 3621 20947 3655
rect 23673 3621 23707 3655
rect 25605 3621 25639 3655
rect 26341 3621 26375 3655
rect 1501 3553 1535 3587
rect 2145 3553 2179 3587
rect 2881 3553 2915 3587
rect 5549 3553 5583 3587
rect 7941 3553 7975 3587
rect 8401 3553 8435 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 10333 3553 10367 3587
rect 10977 3553 11011 3587
rect 11244 3553 11278 3587
rect 12817 3553 12851 3587
rect 13001 3553 13035 3587
rect 13185 3553 13219 3587
rect 15117 3553 15151 3587
rect 15844 3553 15878 3587
rect 17417 3553 17451 3587
rect 18153 3553 18187 3587
rect 18889 3553 18923 3587
rect 19993 3553 20027 3587
rect 20637 3553 20671 3587
rect 20821 3553 20855 3587
rect 21005 3553 21039 3587
rect 21916 3553 21950 3587
rect 23489 3553 23523 3587
rect 23765 3553 23799 3587
rect 23857 3553 23891 3587
rect 26985 3553 27019 3587
rect 15577 3485 15611 3519
rect 21649 3485 21683 3519
rect 7757 3417 7791 3451
rect 12357 3417 12391 3451
rect 25789 3417 25823 3451
rect 26525 3417 26559 3451
rect 1593 3349 1627 3383
rect 3065 3349 3099 3383
rect 8585 3349 8619 3383
rect 10517 3349 10551 3383
rect 13369 3349 13403 3383
rect 16957 3349 16991 3383
rect 18245 3349 18279 3383
rect 20085 3349 20119 3383
rect 21189 3349 21223 3383
rect 23029 3349 23063 3383
rect 24041 3349 24075 3383
rect 4353 3145 4387 3179
rect 5181 3145 5215 3179
rect 13921 3145 13955 3179
rect 18705 3145 18739 3179
rect 21373 3145 21407 3179
rect 24869 3145 24903 3179
rect 1593 3077 1627 3111
rect 12541 3009 12575 3043
rect 19349 3009 19383 3043
rect 23489 3009 23523 3043
rect 1409 2941 1443 2975
rect 2145 2941 2179 2975
rect 2881 2941 2915 2975
rect 3617 2941 3651 2975
rect 4537 2941 4571 2975
rect 4997 2941 5031 2975
rect 6929 2941 6963 2975
rect 8033 2941 8067 2975
rect 8769 2941 8803 2975
rect 9036 2941 9070 2975
rect 10977 2941 11011 2975
rect 12808 2941 12842 2975
rect 14473 2941 14507 2975
rect 15117 2941 15151 2975
rect 15853 2941 15887 2975
rect 16037 2941 16071 2975
rect 16129 2941 16163 2975
rect 16221 2941 16255 2975
rect 17325 2941 17359 2975
rect 21281 2941 21315 2975
rect 22661 2941 22695 2975
rect 23756 2941 23790 2975
rect 25973 2941 26007 2975
rect 26709 2941 26743 2975
rect 11161 2873 11195 2907
rect 17570 2873 17604 2907
rect 19616 2873 19650 2907
rect 26157 2873 26191 2907
rect 10149 2805 10183 2839
rect 14565 2805 14599 2839
rect 16405 2805 16439 2839
rect 20729 2805 20763 2839
rect 22753 2805 22787 2839
rect 26801 2805 26835 2839
rect 5917 2601 5951 2635
rect 12817 2601 12851 2635
rect 16589 2601 16623 2635
rect 19349 2601 19383 2635
rect 22017 2601 22051 2635
rect 23489 2601 23523 2635
rect 25789 2601 25823 2635
rect 27261 2601 27295 2635
rect 4537 2533 4571 2567
rect 10425 2533 10459 2567
rect 12541 2533 12575 2567
rect 16221 2533 16255 2567
rect 16313 2533 16347 2567
rect 17877 2533 17911 2567
rect 18981 2533 19015 2567
rect 20904 2533 20938 2567
rect 23213 2533 23247 2567
rect 25697 2533 25731 2567
rect 26433 2533 26467 2567
rect 1869 2465 1903 2499
rect 2881 2465 2915 2499
rect 4353 2465 4387 2499
rect 4997 2465 5031 2499
rect 5825 2465 5859 2499
rect 7021 2465 7055 2499
rect 7757 2465 7791 2499
rect 8493 2465 8527 2499
rect 9597 2465 9631 2499
rect 11161 2465 11195 2499
rect 12265 2465 12299 2499
rect 12449 2465 12483 2499
rect 12633 2465 12667 2499
rect 13829 2465 13863 2499
rect 15025 2465 15059 2499
rect 16037 2465 16071 2499
rect 16405 2465 16439 2499
rect 17693 2465 17727 2499
rect 18797 2465 18831 2499
rect 19073 2465 19107 2499
rect 19165 2465 19199 2499
rect 20637 2465 20671 2499
rect 22937 2465 22971 2499
rect 23121 2465 23155 2499
rect 23305 2465 23339 2499
rect 24041 2465 24075 2499
rect 27169 2465 27203 2499
rect 11345 2397 11379 2431
rect 3065 2329 3099 2363
rect 5181 2329 5215 2363
rect 7941 2329 7975 2363
rect 8677 2329 8711 2363
rect 10609 2329 10643 2363
rect 15209 2329 15243 2363
rect 26617 2329 26651 2363
rect 1961 2261 1995 2295
rect 7113 2261 7147 2295
rect 13921 2261 13955 2295
rect 24133 2261 24167 2295
<< metal1 >>
rect 15562 29656 15568 29708
rect 15620 29696 15626 29708
rect 27338 29696 27344 29708
rect 15620 29668 27344 29696
rect 15620 29656 15626 29668
rect 27338 29656 27344 29668
rect 27396 29656 27402 29708
rect 9950 29520 9956 29572
rect 10008 29560 10014 29572
rect 20070 29560 20076 29572
rect 10008 29532 20076 29560
rect 10008 29520 10014 29532
rect 20070 29520 20076 29532
rect 20128 29520 20134 29572
rect 15838 29452 15844 29504
rect 15896 29492 15902 29504
rect 21266 29492 21272 29504
rect 15896 29464 21272 29492
rect 15896 29452 15902 29464
rect 21266 29452 21272 29464
rect 21324 29452 21330 29504
rect 1104 29402 28428 29424
rect 1104 29350 5536 29402
rect 5588 29350 5600 29402
rect 5652 29350 5664 29402
rect 5716 29350 5728 29402
rect 5780 29350 14644 29402
rect 14696 29350 14708 29402
rect 14760 29350 14772 29402
rect 14824 29350 14836 29402
rect 14888 29350 23752 29402
rect 23804 29350 23816 29402
rect 23868 29350 23880 29402
rect 23932 29350 23944 29402
rect 23996 29350 28428 29402
rect 1104 29328 28428 29350
rect 3694 29248 3700 29300
rect 3752 29288 3758 29300
rect 4433 29291 4491 29297
rect 4433 29288 4445 29291
rect 3752 29260 4445 29288
rect 3752 29248 3758 29260
rect 4433 29257 4445 29260
rect 4479 29257 4491 29291
rect 4433 29251 4491 29257
rect 5994 29248 6000 29300
rect 6052 29288 6058 29300
rect 7101 29291 7159 29297
rect 7101 29288 7113 29291
rect 6052 29260 7113 29288
rect 6052 29248 6058 29260
rect 7101 29257 7113 29260
rect 7147 29257 7159 29291
rect 7834 29288 7840 29300
rect 7795 29260 7840 29288
rect 7101 29251 7159 29257
rect 7834 29248 7840 29260
rect 7892 29248 7898 29300
rect 10594 29248 10600 29300
rect 10652 29288 10658 29300
rect 10781 29291 10839 29297
rect 10781 29288 10793 29291
rect 10652 29260 10793 29288
rect 10652 29248 10658 29260
rect 10781 29257 10793 29260
rect 10827 29257 10839 29291
rect 10781 29251 10839 29257
rect 12526 29248 12532 29300
rect 12584 29288 12590 29300
rect 13357 29291 13415 29297
rect 13357 29288 13369 29291
rect 12584 29260 13369 29288
rect 12584 29248 12590 29260
rect 13357 29257 13369 29260
rect 13403 29257 13415 29291
rect 13357 29251 13415 29257
rect 15746 29248 15752 29300
rect 15804 29288 15810 29300
rect 16577 29291 16635 29297
rect 16577 29288 16589 29291
rect 15804 29260 16589 29288
rect 15804 29248 15810 29260
rect 16577 29257 16589 29260
rect 16623 29257 16635 29291
rect 16577 29251 16635 29257
rect 17954 29248 17960 29300
rect 18012 29288 18018 29300
rect 18785 29291 18843 29297
rect 18785 29288 18797 29291
rect 18012 29260 18797 29288
rect 18012 29248 18018 29260
rect 18785 29257 18797 29260
rect 18831 29257 18843 29291
rect 18785 29251 18843 29257
rect 20714 29248 20720 29300
rect 20772 29288 20778 29300
rect 20901 29291 20959 29297
rect 20901 29288 20913 29291
rect 20772 29260 20913 29288
rect 20772 29248 20778 29260
rect 20901 29257 20913 29260
rect 20947 29257 20959 29291
rect 20901 29251 20959 29257
rect 21174 29248 21180 29300
rect 21232 29288 21238 29300
rect 21821 29291 21879 29297
rect 21821 29288 21833 29291
rect 21232 29260 21833 29288
rect 21232 29248 21238 29260
rect 21821 29257 21833 29260
rect 21867 29257 21879 29291
rect 21821 29251 21879 29257
rect 22094 29248 22100 29300
rect 22152 29288 22158 29300
rect 23845 29291 23903 29297
rect 23845 29288 23857 29291
rect 22152 29260 23857 29288
rect 22152 29248 22158 29260
rect 23845 29257 23857 29260
rect 23891 29257 23903 29291
rect 23845 29251 23903 29257
rect 24581 29291 24639 29297
rect 24581 29257 24593 29291
rect 24627 29288 24639 29291
rect 28074 29288 28080 29300
rect 24627 29260 28080 29288
rect 24627 29257 24639 29260
rect 24581 29251 24639 29257
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 2406 29180 2412 29232
rect 2464 29220 2470 29232
rect 2685 29223 2743 29229
rect 2685 29220 2697 29223
rect 2464 29192 2697 29220
rect 2464 29180 2470 29192
rect 2685 29189 2697 29192
rect 2731 29189 2743 29223
rect 2685 29183 2743 29189
rect 5813 29223 5871 29229
rect 5813 29189 5825 29223
rect 5859 29220 5871 29223
rect 5902 29220 5908 29232
rect 5859 29192 5908 29220
rect 5859 29189 5871 29192
rect 5813 29183 5871 29189
rect 5902 29180 5908 29192
rect 5960 29180 5966 29232
rect 8665 29223 8723 29229
rect 8665 29189 8677 29223
rect 8711 29220 8723 29223
rect 8754 29220 8760 29232
rect 8711 29192 8760 29220
rect 8711 29189 8723 29192
rect 8665 29183 8723 29189
rect 8754 29180 8760 29192
rect 8812 29180 8818 29232
rect 15933 29223 15991 29229
rect 15933 29189 15945 29223
rect 15979 29220 15991 29223
rect 18874 29220 18880 29232
rect 15979 29192 18880 29220
rect 15979 29189 15991 29192
rect 15933 29183 15991 29189
rect 18874 29180 18880 29192
rect 18932 29180 18938 29232
rect 19794 29180 19800 29232
rect 19852 29220 19858 29232
rect 23201 29223 23259 29229
rect 23201 29220 23213 29223
rect 19852 29192 23213 29220
rect 19852 29180 19858 29192
rect 23201 29189 23213 29192
rect 23247 29189 23259 29223
rect 23201 29183 23259 29189
rect 25869 29223 25927 29229
rect 25869 29189 25881 29223
rect 25915 29220 25927 29223
rect 27614 29220 27620 29232
rect 25915 29192 27620 29220
rect 25915 29189 25927 29192
rect 25869 29183 25927 29189
rect 27614 29180 27620 29192
rect 27672 29180 27678 29232
rect 2958 29112 2964 29164
rect 3016 29152 3022 29164
rect 3016 29124 17816 29152
rect 3016 29112 3022 29124
rect 1854 29084 1860 29096
rect 1815 29056 1860 29084
rect 1854 29044 1860 29056
rect 1912 29044 1918 29096
rect 1946 29044 1952 29096
rect 2004 29084 2010 29096
rect 2501 29087 2559 29093
rect 2501 29084 2513 29087
rect 2004 29056 2513 29084
rect 2004 29044 2010 29056
rect 2501 29053 2513 29056
rect 2547 29053 2559 29087
rect 2501 29047 2559 29053
rect 7009 29087 7067 29093
rect 7009 29053 7021 29087
rect 7055 29084 7067 29087
rect 9950 29084 9956 29096
rect 7055 29056 9812 29084
rect 9911 29056 9956 29084
rect 7055 29053 7067 29056
rect 7009 29047 7067 29053
rect 2041 29019 2099 29025
rect 2041 28985 2053 29019
rect 2087 29016 2099 29019
rect 2222 29016 2228 29028
rect 2087 28988 2228 29016
rect 2087 28985 2099 28988
rect 2041 28979 2099 28985
rect 2222 28976 2228 28988
rect 2280 28976 2286 29028
rect 4341 29019 4399 29025
rect 4341 28985 4353 29019
rect 4387 29016 4399 29019
rect 5350 29016 5356 29028
rect 4387 28988 5356 29016
rect 4387 28985 4399 28988
rect 4341 28979 4399 28985
rect 5350 28976 5356 28988
rect 5408 28976 5414 29028
rect 5626 29016 5632 29028
rect 5587 28988 5632 29016
rect 5626 28976 5632 28988
rect 5684 28976 5690 29028
rect 7742 29016 7748 29028
rect 7703 28988 7748 29016
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 8481 29019 8539 29025
rect 8481 28985 8493 29019
rect 8527 28985 8539 29019
rect 9784 29016 9812 29056
rect 9950 29044 9956 29056
rect 10008 29044 10014 29096
rect 10137 29087 10195 29093
rect 10137 29053 10149 29087
rect 10183 29084 10195 29087
rect 10962 29084 10968 29096
rect 10183 29056 10968 29084
rect 10183 29053 10195 29056
rect 10137 29047 10195 29053
rect 10962 29044 10968 29056
rect 11020 29044 11026 29096
rect 12434 29044 12440 29096
rect 12492 29084 12498 29096
rect 12529 29087 12587 29093
rect 12529 29084 12541 29087
rect 12492 29056 12541 29084
rect 12492 29044 12498 29056
rect 12529 29053 12541 29056
rect 12575 29053 12587 29087
rect 12529 29047 12587 29053
rect 12894 29044 12900 29096
rect 12952 29084 12958 29096
rect 13265 29087 13323 29093
rect 13265 29084 13277 29087
rect 12952 29056 13277 29084
rect 12952 29044 12958 29056
rect 13265 29053 13277 29056
rect 13311 29053 13323 29087
rect 15010 29084 15016 29096
rect 14971 29056 15016 29084
rect 13265 29047 13323 29053
rect 15010 29044 15016 29056
rect 15068 29044 15074 29096
rect 15197 29087 15255 29093
rect 15197 29053 15209 29087
rect 15243 29084 15255 29087
rect 16298 29084 16304 29096
rect 15243 29056 16304 29084
rect 15243 29053 15255 29056
rect 15197 29047 15255 29053
rect 16298 29044 16304 29056
rect 16356 29044 16362 29096
rect 16393 29087 16451 29093
rect 16393 29053 16405 29087
rect 16439 29084 16451 29087
rect 17034 29084 17040 29096
rect 16439 29056 17040 29084
rect 16439 29053 16451 29056
rect 16393 29047 16451 29053
rect 17034 29044 17040 29056
rect 17092 29044 17098 29096
rect 17589 29087 17647 29093
rect 17589 29053 17601 29087
rect 17635 29084 17647 29087
rect 17678 29084 17684 29096
rect 17635 29056 17684 29084
rect 17635 29053 17647 29056
rect 17589 29047 17647 29053
rect 17678 29044 17684 29056
rect 17736 29044 17742 29096
rect 17788 29093 17816 29124
rect 18800 29124 19656 29152
rect 18046 29093 18052 29096
rect 17773 29087 17831 29093
rect 17773 29053 17785 29087
rect 17819 29053 17831 29087
rect 17773 29047 17831 29053
rect 18003 29087 18052 29093
rect 18003 29053 18015 29087
rect 18049 29053 18052 29087
rect 18003 29047 18052 29053
rect 18046 29044 18052 29047
rect 18104 29044 18110 29096
rect 18693 29087 18751 29093
rect 18693 29053 18705 29087
rect 18739 29084 18751 29087
rect 18800 29084 18828 29124
rect 18739 29056 18828 29084
rect 19628 29084 19656 29124
rect 19702 29112 19708 29164
rect 19760 29152 19766 29164
rect 27338 29152 27344 29164
rect 19760 29124 23060 29152
rect 27299 29124 27344 29152
rect 19760 29112 19766 29124
rect 19628 29056 20944 29084
rect 18739 29053 18751 29056
rect 18693 29047 18751 29053
rect 9858 29016 9864 29028
rect 9784 28988 9864 29016
rect 8481 28979 8539 28985
rect 6914 28908 6920 28960
rect 6972 28948 6978 28960
rect 8294 28948 8300 28960
rect 6972 28920 8300 28948
rect 6972 28908 6978 28920
rect 8294 28908 8300 28920
rect 8352 28908 8358 28960
rect 8496 28948 8524 28979
rect 9858 28976 9864 28988
rect 9916 28976 9922 29028
rect 10686 29016 10692 29028
rect 9968 28988 10180 29016
rect 10647 28988 10692 29016
rect 9490 28948 9496 28960
rect 8496 28920 9496 28948
rect 9490 28908 9496 28920
rect 9548 28948 9554 28960
rect 9968 28948 9996 28988
rect 9548 28920 9996 28948
rect 10152 28948 10180 28988
rect 10686 28976 10692 28988
rect 10744 28976 10750 29028
rect 12713 29019 12771 29025
rect 12713 28985 12725 29019
rect 12759 29016 12771 29019
rect 12802 29016 12808 29028
rect 12759 28988 12808 29016
rect 12759 28985 12771 28988
rect 12713 28979 12771 28985
rect 12802 28976 12808 28988
rect 12860 28976 12866 29028
rect 15749 29019 15807 29025
rect 15749 28985 15761 29019
rect 15795 29016 15807 29019
rect 15838 29016 15844 29028
rect 15795 28988 15844 29016
rect 15795 28985 15807 28988
rect 15749 28979 15807 28985
rect 15838 28976 15844 28988
rect 15896 28976 15902 29028
rect 17861 29019 17919 29025
rect 17861 28985 17873 29019
rect 17907 28985 17919 29019
rect 18782 29016 18788 29028
rect 17861 28979 17919 28985
rect 17972 28988 18788 29016
rect 16022 28948 16028 28960
rect 10152 28920 16028 28948
rect 9548 28908 9554 28920
rect 16022 28908 16028 28920
rect 16080 28908 16086 28960
rect 17880 28948 17908 28979
rect 17972 28948 18000 28988
rect 18782 28976 18788 28988
rect 18840 28976 18846 29028
rect 20809 29019 20867 29025
rect 20809 28985 20821 29019
rect 20855 28985 20867 29019
rect 20916 29016 20944 29056
rect 21634 29044 21640 29096
rect 21692 29084 21698 29096
rect 23032 29093 23060 29124
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 21729 29087 21787 29093
rect 21729 29084 21741 29087
rect 21692 29056 21741 29084
rect 21692 29044 21698 29056
rect 21729 29053 21741 29056
rect 21775 29053 21787 29087
rect 21729 29047 21787 29053
rect 23017 29087 23075 29093
rect 23017 29053 23029 29087
rect 23063 29053 23075 29087
rect 23017 29047 23075 29053
rect 24489 29087 24547 29093
rect 24489 29053 24501 29087
rect 24535 29084 24547 29087
rect 25958 29084 25964 29096
rect 24535 29056 25964 29084
rect 24535 29053 24547 29056
rect 24489 29047 24547 29053
rect 25958 29044 25964 29056
rect 26016 29044 26022 29096
rect 26142 29044 26148 29096
rect 26200 29084 26206 29096
rect 26421 29087 26479 29093
rect 26421 29084 26433 29087
rect 26200 29056 26433 29084
rect 26200 29044 26206 29056
rect 26421 29053 26433 29056
rect 26467 29053 26479 29087
rect 27154 29084 27160 29096
rect 27115 29056 27160 29084
rect 26421 29047 26479 29053
rect 27154 29044 27160 29056
rect 27212 29044 27218 29096
rect 23750 29016 23756 29028
rect 20916 28988 23612 29016
rect 23711 28988 23756 29016
rect 20809 28979 20867 28985
rect 18138 28948 18144 28960
rect 17880 28920 18000 28948
rect 18099 28920 18144 28948
rect 18138 28908 18144 28920
rect 18196 28908 18202 28960
rect 20824 28948 20852 28979
rect 20990 28948 20996 28960
rect 20824 28920 20996 28948
rect 20990 28908 20996 28920
rect 21048 28908 21054 28960
rect 23584 28948 23612 28988
rect 23750 28976 23756 28988
rect 23808 28976 23814 29028
rect 25590 28976 25596 29028
rect 25648 29016 25654 29028
rect 25685 29019 25743 29025
rect 25685 29016 25697 29019
rect 25648 28988 25697 29016
rect 25648 28976 25654 28988
rect 25685 28985 25697 28988
rect 25731 28985 25743 29019
rect 25685 28979 25743 28985
rect 26605 29019 26663 29025
rect 26605 28985 26617 29019
rect 26651 29016 26663 29019
rect 26786 29016 26792 29028
rect 26651 28988 26792 29016
rect 26651 28985 26663 28988
rect 26605 28979 26663 28985
rect 26786 28976 26792 28988
rect 26844 28976 26850 29028
rect 24578 28948 24584 28960
rect 23584 28920 24584 28948
rect 24578 28908 24584 28920
rect 24636 28908 24642 28960
rect 1104 28858 28428 28880
rect 1104 28806 10090 28858
rect 10142 28806 10154 28858
rect 10206 28806 10218 28858
rect 10270 28806 10282 28858
rect 10334 28806 19198 28858
rect 19250 28806 19262 28858
rect 19314 28806 19326 28858
rect 19378 28806 19390 28858
rect 19442 28806 28428 28858
rect 1104 28784 28428 28806
rect 474 28704 480 28756
rect 532 28744 538 28756
rect 1949 28747 2007 28753
rect 1949 28744 1961 28747
rect 532 28716 1961 28744
rect 532 28704 538 28716
rect 1949 28713 1961 28716
rect 1995 28713 2007 28747
rect 1949 28707 2007 28713
rect 2314 28704 2320 28756
rect 2372 28744 2378 28756
rect 3053 28747 3111 28753
rect 3053 28744 3065 28747
rect 2372 28716 3065 28744
rect 2372 28704 2378 28716
rect 3053 28713 3065 28716
rect 3099 28713 3111 28747
rect 3053 28707 3111 28713
rect 5626 28704 5632 28756
rect 5684 28744 5690 28756
rect 5684 28716 15976 28744
rect 5684 28704 5690 28716
rect 1762 28568 1768 28620
rect 1820 28608 1826 28620
rect 1857 28611 1915 28617
rect 1857 28608 1869 28611
rect 1820 28580 1869 28608
rect 1820 28568 1826 28580
rect 1857 28577 1869 28580
rect 1903 28577 1915 28611
rect 1857 28571 1915 28577
rect 2961 28611 3019 28617
rect 2961 28577 2973 28611
rect 3007 28608 3019 28611
rect 3418 28608 3424 28620
rect 3007 28580 3424 28608
rect 3007 28577 3019 28580
rect 2961 28571 3019 28577
rect 3418 28568 3424 28580
rect 3476 28568 3482 28620
rect 4154 28568 4160 28620
rect 4212 28608 4218 28620
rect 4249 28611 4307 28617
rect 4249 28608 4261 28611
rect 4212 28580 4261 28608
rect 4212 28568 4218 28580
rect 4249 28577 4261 28580
rect 4295 28577 4307 28611
rect 5074 28608 5080 28620
rect 5035 28580 5080 28608
rect 4249 28571 4307 28577
rect 5074 28568 5080 28580
rect 5132 28568 5138 28620
rect 6196 28617 6224 28716
rect 7466 28676 7472 28688
rect 7427 28648 7472 28676
rect 7466 28636 7472 28648
rect 7524 28636 7530 28688
rect 9674 28636 9680 28688
rect 9732 28676 9738 28688
rect 9732 28648 10916 28676
rect 9732 28636 9738 28648
rect 6181 28611 6239 28617
rect 6181 28577 6193 28611
rect 6227 28577 6239 28611
rect 6181 28571 6239 28577
rect 7098 28568 7104 28620
rect 7156 28608 7162 28620
rect 7285 28611 7343 28617
rect 7285 28608 7297 28611
rect 7156 28580 7297 28608
rect 7156 28568 7162 28580
rect 7285 28577 7297 28580
rect 7331 28577 7343 28611
rect 7558 28608 7564 28620
rect 7519 28580 7564 28608
rect 7285 28571 7343 28577
rect 7558 28568 7564 28580
rect 7616 28568 7622 28620
rect 7699 28611 7757 28617
rect 7699 28577 7711 28611
rect 7745 28608 7757 28611
rect 7834 28608 7840 28620
rect 7745 28580 7840 28608
rect 7745 28577 7757 28580
rect 7699 28571 7757 28577
rect 7834 28568 7840 28580
rect 7892 28568 7898 28620
rect 8294 28608 8300 28620
rect 8255 28580 8300 28608
rect 8294 28568 8300 28580
rect 8352 28568 8358 28620
rect 9490 28608 9496 28620
rect 9451 28580 9496 28608
rect 9490 28568 9496 28580
rect 9548 28568 9554 28620
rect 10502 28617 10508 28620
rect 10496 28571 10508 28617
rect 10560 28608 10566 28620
rect 10888 28608 10916 28648
rect 11054 28636 11060 28688
rect 11112 28676 11118 28688
rect 15948 28676 15976 28716
rect 16022 28704 16028 28756
rect 16080 28744 16086 28756
rect 16117 28747 16175 28753
rect 16117 28744 16129 28747
rect 16080 28716 16129 28744
rect 16080 28704 16086 28716
rect 16117 28713 16129 28716
rect 16163 28744 16175 28747
rect 16390 28744 16396 28756
rect 16163 28716 16396 28744
rect 16163 28713 16175 28716
rect 16117 28707 16175 28713
rect 16390 28704 16396 28716
rect 16448 28704 16454 28756
rect 17586 28676 17592 28688
rect 11112 28648 12434 28676
rect 15948 28648 17592 28676
rect 11112 28636 11118 28648
rect 12069 28611 12127 28617
rect 12069 28608 12081 28611
rect 10560 28580 10596 28608
rect 10888 28580 12081 28608
rect 10502 28568 10508 28571
rect 10560 28568 10566 28580
rect 12069 28577 12081 28580
rect 12115 28577 12127 28611
rect 12406 28608 12434 28648
rect 17586 28636 17592 28648
rect 17644 28636 17650 28688
rect 20254 28636 20260 28688
rect 20312 28676 20318 28688
rect 24305 28679 24363 28685
rect 20312 28648 22094 28676
rect 20312 28636 20318 28648
rect 12897 28611 12955 28617
rect 12897 28608 12909 28611
rect 12406 28580 12909 28608
rect 12069 28571 12127 28577
rect 12897 28577 12909 28580
rect 12943 28577 12955 28611
rect 13354 28608 13360 28620
rect 13315 28580 13360 28608
rect 12897 28571 12955 28577
rect 13354 28568 13360 28580
rect 13412 28568 13418 28620
rect 15004 28611 15062 28617
rect 15004 28577 15016 28611
rect 15050 28608 15062 28611
rect 16022 28608 16028 28620
rect 15050 28580 16028 28608
rect 15050 28577 15062 28580
rect 15004 28571 15062 28577
rect 16022 28568 16028 28580
rect 16080 28568 16086 28620
rect 16114 28568 16120 28620
rect 16172 28608 16178 28620
rect 16577 28611 16635 28617
rect 16577 28608 16589 28611
rect 16172 28580 16589 28608
rect 16172 28568 16178 28580
rect 16577 28577 16589 28580
rect 16623 28577 16635 28611
rect 16577 28571 16635 28577
rect 17764 28611 17822 28617
rect 17764 28577 17776 28611
rect 17810 28608 17822 28611
rect 18046 28608 18052 28620
rect 17810 28580 18052 28608
rect 17810 28577 17822 28580
rect 17764 28571 17822 28577
rect 18046 28568 18052 28580
rect 18104 28568 18110 28620
rect 20070 28608 20076 28620
rect 20031 28580 20076 28608
rect 20070 28568 20076 28580
rect 20128 28568 20134 28620
rect 20809 28611 20867 28617
rect 20809 28577 20821 28611
rect 20855 28608 20867 28611
rect 20990 28608 20996 28620
rect 20855 28580 20996 28608
rect 20855 28577 20867 28580
rect 20809 28571 20867 28577
rect 20990 28568 20996 28580
rect 21048 28568 21054 28620
rect 21545 28611 21603 28617
rect 21545 28577 21557 28611
rect 21591 28577 21603 28611
rect 22066 28608 22094 28648
rect 24305 28645 24317 28679
rect 24351 28676 24363 28679
rect 24394 28676 24400 28688
rect 24351 28648 24400 28676
rect 24351 28645 24363 28648
rect 24305 28639 24363 28645
rect 24394 28636 24400 28648
rect 24452 28636 24458 28688
rect 25777 28679 25835 28685
rect 25777 28645 25789 28679
rect 25823 28676 25835 28679
rect 28994 28676 29000 28688
rect 25823 28648 29000 28676
rect 25823 28645 25835 28648
rect 25777 28639 25835 28645
rect 28994 28636 29000 28648
rect 29052 28636 29058 28688
rect 22281 28611 22339 28617
rect 22281 28608 22293 28611
rect 22066 28580 22293 28608
rect 21545 28571 21603 28577
rect 22281 28577 22293 28580
rect 22327 28577 22339 28611
rect 22281 28571 22339 28577
rect 23385 28611 23443 28617
rect 23385 28577 23397 28611
rect 23431 28608 23443 28611
rect 23474 28608 23480 28620
rect 23431 28580 23480 28608
rect 23431 28577 23443 28580
rect 23385 28571 23443 28577
rect 8570 28500 8576 28552
rect 8628 28540 8634 28552
rect 9950 28540 9956 28552
rect 8628 28512 9956 28540
rect 8628 28500 8634 28512
rect 9950 28500 9956 28512
rect 10008 28500 10014 28552
rect 10226 28540 10232 28552
rect 10187 28512 10232 28540
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 14458 28500 14464 28552
rect 14516 28540 14522 28552
rect 14737 28543 14795 28549
rect 14737 28540 14749 28543
rect 14516 28512 14749 28540
rect 14516 28500 14522 28512
rect 14737 28509 14749 28512
rect 14783 28509 14795 28543
rect 14737 28503 14795 28509
rect 17218 28500 17224 28552
rect 17276 28540 17282 28552
rect 17497 28543 17555 28549
rect 17497 28540 17509 28543
rect 17276 28512 17509 28540
rect 17276 28500 17282 28512
rect 17497 28509 17509 28512
rect 17543 28509 17555 28543
rect 17497 28503 17555 28509
rect 20898 28500 20904 28552
rect 20956 28540 20962 28552
rect 21560 28540 21588 28571
rect 23474 28568 23480 28580
rect 23532 28568 23538 28620
rect 24121 28611 24179 28617
rect 24121 28577 24133 28611
rect 24167 28608 24179 28611
rect 24210 28608 24216 28620
rect 24167 28580 24216 28608
rect 24167 28577 24179 28580
rect 24121 28571 24179 28577
rect 24210 28568 24216 28580
rect 24268 28568 24274 28620
rect 25038 28568 25044 28620
rect 25096 28608 25102 28620
rect 25593 28611 25651 28617
rect 25593 28608 25605 28611
rect 25096 28580 25605 28608
rect 25096 28568 25102 28580
rect 25593 28577 25605 28580
rect 25639 28577 25651 28611
rect 25593 28571 25651 28577
rect 26329 28611 26387 28617
rect 26329 28577 26341 28611
rect 26375 28608 26387 28611
rect 26418 28608 26424 28620
rect 26375 28580 26424 28608
rect 26375 28577 26387 28580
rect 26329 28571 26387 28577
rect 23750 28540 23756 28552
rect 20956 28512 23756 28540
rect 20956 28500 20962 28512
rect 23750 28500 23756 28512
rect 23808 28500 23814 28552
rect 25608 28540 25636 28571
rect 26418 28568 26424 28580
rect 26476 28568 26482 28620
rect 26973 28611 27031 28617
rect 26973 28577 26985 28611
rect 27019 28577 27031 28611
rect 26973 28571 27031 28577
rect 26988 28540 27016 28571
rect 25608 28512 27016 28540
rect 5261 28475 5319 28481
rect 5261 28441 5273 28475
rect 5307 28472 5319 28475
rect 9858 28472 9864 28484
rect 5307 28444 9864 28472
rect 5307 28441 5319 28444
rect 5261 28435 5319 28441
rect 9858 28432 9864 28444
rect 9916 28432 9922 28484
rect 17402 28472 17408 28484
rect 16040 28444 17408 28472
rect 4433 28407 4491 28413
rect 4433 28373 4445 28407
rect 4479 28404 4491 28407
rect 4982 28404 4988 28416
rect 4479 28376 4988 28404
rect 4479 28373 4491 28376
rect 4433 28367 4491 28373
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 7466 28364 7472 28416
rect 7524 28404 7530 28416
rect 7837 28407 7895 28413
rect 7837 28404 7849 28407
rect 7524 28376 7849 28404
rect 7524 28364 7530 28376
rect 7837 28373 7849 28376
rect 7883 28373 7895 28407
rect 7837 28367 7895 28373
rect 8481 28407 8539 28413
rect 8481 28373 8493 28407
rect 8527 28404 8539 28407
rect 10410 28404 10416 28416
rect 8527 28376 10416 28404
rect 8527 28373 8539 28376
rect 8481 28367 8539 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 11146 28364 11152 28416
rect 11204 28404 11210 28416
rect 11609 28407 11667 28413
rect 11609 28404 11621 28407
rect 11204 28376 11621 28404
rect 11204 28364 11210 28376
rect 11609 28373 11621 28376
rect 11655 28373 11667 28407
rect 11609 28367 11667 28373
rect 12713 28407 12771 28413
rect 12713 28373 12725 28407
rect 12759 28404 12771 28407
rect 16040 28404 16068 28444
rect 17402 28432 17408 28444
rect 17460 28432 17466 28484
rect 22465 28475 22523 28481
rect 22465 28472 22477 28475
rect 18432 28444 22477 28472
rect 12759 28376 16068 28404
rect 12759 28373 12771 28376
rect 12713 28367 12771 28373
rect 17494 28364 17500 28416
rect 17552 28404 17558 28416
rect 18432 28404 18460 28444
rect 22465 28441 22477 28444
rect 22511 28441 22523 28475
rect 22465 28435 22523 28441
rect 18874 28404 18880 28416
rect 17552 28376 18460 28404
rect 18835 28376 18880 28404
rect 17552 28364 17558 28376
rect 18874 28364 18880 28376
rect 18932 28364 18938 28416
rect 22646 28364 22652 28416
rect 22704 28404 22710 28416
rect 23569 28407 23627 28413
rect 23569 28404 23581 28407
rect 22704 28376 23581 28404
rect 22704 28364 22710 28376
rect 23569 28373 23581 28376
rect 23615 28373 23627 28407
rect 23569 28367 23627 28373
rect 26142 28364 26148 28416
rect 26200 28404 26206 28416
rect 26421 28407 26479 28413
rect 26421 28404 26433 28407
rect 26200 28376 26433 28404
rect 26200 28364 26206 28376
rect 26421 28373 26433 28376
rect 26467 28373 26479 28407
rect 26421 28367 26479 28373
rect 1104 28314 28428 28336
rect 1104 28262 5536 28314
rect 5588 28262 5600 28314
rect 5652 28262 5664 28314
rect 5716 28262 5728 28314
rect 5780 28262 14644 28314
rect 14696 28262 14708 28314
rect 14760 28262 14772 28314
rect 14824 28262 14836 28314
rect 14888 28262 23752 28314
rect 23804 28262 23816 28314
rect 23868 28262 23880 28314
rect 23932 28262 23944 28314
rect 23996 28262 28428 28314
rect 1104 28240 28428 28262
rect 2317 28203 2375 28209
rect 2317 28169 2329 28203
rect 2363 28200 2375 28203
rect 2363 28172 20484 28200
rect 2363 28169 2375 28172
rect 2317 28163 2375 28169
rect 2774 28092 2780 28144
rect 2832 28092 2838 28144
rect 2958 28132 2964 28144
rect 2919 28104 2964 28132
rect 2958 28092 2964 28104
rect 3016 28092 3022 28144
rect 10410 28092 10416 28144
rect 10468 28132 10474 28144
rect 12986 28132 12992 28144
rect 10468 28104 12992 28132
rect 10468 28092 10474 28104
rect 12986 28092 12992 28104
rect 13044 28092 13050 28144
rect 18782 28092 18788 28144
rect 18840 28132 18846 28144
rect 18877 28135 18935 28141
rect 18877 28132 18889 28135
rect 18840 28104 18889 28132
rect 18840 28092 18846 28104
rect 18877 28101 18889 28104
rect 18923 28101 18935 28135
rect 18877 28095 18935 28101
rect 2792 28064 2820 28092
rect 10226 28064 10232 28076
rect 2792 28036 3648 28064
rect 1394 27996 1400 28008
rect 1355 27968 1400 27996
rect 1394 27956 1400 27968
rect 1452 27956 1458 28008
rect 2130 27996 2136 28008
rect 2091 27968 2136 27996
rect 2130 27956 2136 27968
rect 2188 27956 2194 28008
rect 2774 27956 2780 28008
rect 2832 27996 2838 28008
rect 3620 28005 3648 28036
rect 9692 28036 10232 28064
rect 3605 27999 3663 28005
rect 2832 27968 2877 27996
rect 2832 27956 2838 27968
rect 3605 27965 3617 27999
rect 3651 27965 3663 27999
rect 3605 27959 3663 27965
rect 6825 27999 6883 28005
rect 6825 27965 6837 27999
rect 6871 27965 6883 27999
rect 6825 27959 6883 27965
rect 7092 27999 7150 28005
rect 7092 27965 7104 27999
rect 7138 27996 7150 27999
rect 7466 27996 7472 28008
rect 7138 27968 7472 27996
rect 7138 27965 7150 27968
rect 7092 27959 7150 27965
rect 6840 27928 6868 27959
rect 7466 27956 7472 27968
rect 7524 27956 7530 28008
rect 8665 27999 8723 28005
rect 8665 27965 8677 27999
rect 8711 27996 8723 27999
rect 9490 27996 9496 28008
rect 8711 27968 9496 27996
rect 8711 27965 8723 27968
rect 8665 27959 8723 27965
rect 8680 27928 8708 27959
rect 9490 27956 9496 27968
rect 9548 27996 9554 28008
rect 9692 27996 9720 28036
rect 10226 28024 10232 28036
rect 10284 28024 10290 28076
rect 9548 27968 9720 27996
rect 10505 27999 10563 28005
rect 9548 27956 9554 27968
rect 10505 27965 10517 27999
rect 10551 27996 10563 27999
rect 10686 27996 10692 28008
rect 10551 27968 10692 27996
rect 10551 27965 10563 27968
rect 10505 27959 10563 27965
rect 6840 27900 8708 27928
rect 8754 27888 8760 27940
rect 8812 27928 8818 27940
rect 8910 27931 8968 27937
rect 8910 27928 8922 27931
rect 8812 27900 8922 27928
rect 8812 27888 8818 27900
rect 8910 27897 8922 27900
rect 8956 27897 8968 27931
rect 8910 27891 8968 27897
rect 9674 27888 9680 27940
rect 9732 27928 9738 27940
rect 10520 27928 10548 27959
rect 10686 27956 10692 27968
rect 10744 27956 10750 28008
rect 11514 27956 11520 28008
rect 11572 27996 11578 28008
rect 12069 27999 12127 28005
rect 12069 27996 12081 27999
rect 11572 27968 12081 27996
rect 11572 27956 11578 27968
rect 12069 27965 12081 27968
rect 12115 27965 12127 27999
rect 12069 27959 12127 27965
rect 13909 27999 13967 28005
rect 13909 27965 13921 27999
rect 13955 27965 13967 27999
rect 14366 27996 14372 28008
rect 14327 27968 14372 27996
rect 13909 27959 13967 27965
rect 9732 27900 10548 27928
rect 13924 27928 13952 27959
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 15194 27996 15200 28008
rect 14476 27968 15200 27996
rect 14476 27928 14504 27968
rect 15194 27956 15200 27968
rect 15252 27956 15258 28008
rect 17218 27956 17224 28008
rect 17276 27996 17282 28008
rect 17497 27999 17555 28005
rect 17497 27996 17509 27999
rect 17276 27968 17509 27996
rect 17276 27956 17282 27968
rect 17497 27965 17509 27968
rect 17543 27965 17555 27999
rect 17497 27959 17555 27965
rect 17764 27999 17822 28005
rect 17764 27965 17776 27999
rect 17810 27996 17822 27999
rect 18138 27996 18144 28008
rect 17810 27968 18144 27996
rect 17810 27965 17822 27968
rect 17764 27959 17822 27965
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 19337 27999 19395 28005
rect 19337 27965 19349 27999
rect 19383 27996 19395 27999
rect 19702 27996 19708 28008
rect 19383 27968 19708 27996
rect 19383 27965 19395 27968
rect 19337 27959 19395 27965
rect 19702 27956 19708 27968
rect 19760 27956 19766 28008
rect 20456 28005 20484 28172
rect 21726 28064 21732 28076
rect 20548 28036 21732 28064
rect 20548 28005 20576 28036
rect 21726 28024 21732 28036
rect 21784 28024 21790 28076
rect 20257 27999 20315 28005
rect 20257 27965 20269 27999
rect 20303 27965 20315 27999
rect 20257 27959 20315 27965
rect 20441 27999 20499 28005
rect 20441 27965 20453 27999
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 20533 27999 20591 28005
rect 20533 27965 20545 27999
rect 20579 27965 20591 27999
rect 20533 27959 20591 27965
rect 20625 27999 20683 28005
rect 20625 27965 20637 27999
rect 20671 27965 20683 27999
rect 21266 27996 21272 28008
rect 21179 27968 21272 27996
rect 20625 27959 20683 27965
rect 13924 27900 14504 27928
rect 14636 27931 14694 27937
rect 9732 27888 9738 27900
rect 14636 27897 14648 27931
rect 14682 27928 14694 27931
rect 15286 27928 15292 27940
rect 14682 27900 15292 27928
rect 14682 27897 14694 27900
rect 14636 27891 14694 27897
rect 15286 27888 15292 27900
rect 15344 27888 15350 27940
rect 17678 27888 17684 27940
rect 17736 27928 17742 27940
rect 20272 27928 20300 27959
rect 17736 27900 20300 27928
rect 17736 27888 17742 27900
rect 3421 27863 3479 27869
rect 3421 27829 3433 27863
rect 3467 27860 3479 27863
rect 4430 27860 4436 27872
rect 3467 27832 4436 27860
rect 3467 27829 3479 27832
rect 3421 27823 3479 27829
rect 4430 27820 4436 27832
rect 4488 27820 4494 27872
rect 6638 27820 6644 27872
rect 6696 27860 6702 27872
rect 7558 27860 7564 27872
rect 6696 27832 7564 27860
rect 6696 27820 6702 27832
rect 7558 27820 7564 27832
rect 7616 27860 7622 27872
rect 8205 27863 8263 27869
rect 8205 27860 8217 27863
rect 7616 27832 8217 27860
rect 7616 27820 7622 27832
rect 8205 27829 8217 27832
rect 8251 27829 8263 27863
rect 8205 27823 8263 27829
rect 9766 27820 9772 27872
rect 9824 27860 9830 27872
rect 10045 27863 10103 27869
rect 10045 27860 10057 27863
rect 9824 27832 10057 27860
rect 9824 27820 9830 27832
rect 10045 27829 10057 27832
rect 10091 27829 10103 27863
rect 10045 27823 10103 27829
rect 10410 27820 10416 27872
rect 10468 27860 10474 27872
rect 12253 27863 12311 27869
rect 12253 27860 12265 27863
rect 10468 27832 12265 27860
rect 10468 27820 10474 27832
rect 12253 27829 12265 27832
rect 12299 27829 12311 27863
rect 12253 27823 12311 27829
rect 13078 27820 13084 27872
rect 13136 27860 13142 27872
rect 13725 27863 13783 27869
rect 13725 27860 13737 27863
rect 13136 27832 13737 27860
rect 13136 27820 13142 27832
rect 13725 27829 13737 27832
rect 13771 27829 13783 27863
rect 13725 27823 13783 27829
rect 15378 27820 15384 27872
rect 15436 27860 15442 27872
rect 15749 27863 15807 27869
rect 15749 27860 15761 27863
rect 15436 27832 15761 27860
rect 15436 27820 15442 27832
rect 15749 27829 15761 27832
rect 15795 27860 15807 27863
rect 16114 27860 16120 27872
rect 15795 27832 16120 27860
rect 15795 27829 15807 27832
rect 15749 27823 15807 27829
rect 16114 27820 16120 27832
rect 16172 27820 16178 27872
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 20640 27860 20668 27959
rect 21266 27956 21272 27968
rect 21324 27996 21330 28008
rect 21634 27996 21640 28008
rect 21324 27968 21640 27996
rect 21324 27956 21330 27968
rect 21634 27956 21640 27968
rect 21692 27956 21698 28008
rect 22554 27996 22560 28008
rect 22515 27968 22560 27996
rect 22554 27956 22560 27968
rect 22612 27956 22618 28008
rect 23937 27999 23995 28005
rect 23937 27965 23949 27999
rect 23983 27996 23995 27999
rect 24118 27996 24124 28008
rect 23983 27968 24124 27996
rect 23983 27965 23995 27968
rect 23937 27959 23995 27965
rect 24118 27956 24124 27968
rect 24176 27956 24182 28008
rect 24578 27996 24584 28008
rect 24539 27968 24584 27996
rect 24578 27956 24584 27968
rect 24636 27956 24642 28008
rect 25314 27996 25320 28008
rect 25275 27968 25320 27996
rect 25314 27956 25320 27968
rect 25372 27956 25378 28008
rect 25958 27996 25964 28008
rect 25919 27968 25964 27996
rect 25958 27956 25964 27968
rect 26016 27956 26022 28008
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 26697 27999 26755 28005
rect 26697 27996 26709 27999
rect 26292 27968 26709 27996
rect 26292 27956 26298 27968
rect 26697 27965 26709 27968
rect 26743 27965 26755 27999
rect 26697 27959 26755 27965
rect 20806 27860 20812 27872
rect 18012 27832 20668 27860
rect 20767 27832 20812 27860
rect 18012 27820 18018 27832
rect 20806 27820 20812 27832
rect 20864 27820 20870 27872
rect 22370 27820 22376 27872
rect 22428 27860 22434 27872
rect 22741 27863 22799 27869
rect 22741 27860 22753 27863
rect 22428 27832 22753 27860
rect 22428 27820 22434 27832
rect 22741 27829 22753 27832
rect 22787 27829 22799 27863
rect 22741 27823 22799 27829
rect 24121 27863 24179 27869
rect 24121 27829 24133 27863
rect 24167 27860 24179 27863
rect 24670 27860 24676 27872
rect 24167 27832 24676 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 24670 27820 24676 27832
rect 24728 27820 24734 27872
rect 1104 27770 28428 27792
rect 1104 27718 10090 27770
rect 10142 27718 10154 27770
rect 10206 27718 10218 27770
rect 10270 27718 10282 27770
rect 10334 27718 19198 27770
rect 19250 27718 19262 27770
rect 19314 27718 19326 27770
rect 19378 27718 19390 27770
rect 19442 27718 28428 27770
rect 1104 27696 28428 27718
rect 10502 27616 10508 27668
rect 10560 27656 10566 27668
rect 10689 27659 10747 27665
rect 10689 27656 10701 27659
rect 10560 27628 10701 27656
rect 10560 27616 10566 27628
rect 10689 27625 10701 27628
rect 10735 27625 10747 27659
rect 12250 27656 12256 27668
rect 10689 27619 10747 27625
rect 10888 27628 12256 27656
rect 934 27548 940 27600
rect 992 27588 998 27600
rect 2774 27588 2780 27600
rect 992 27560 2780 27588
rect 992 27548 998 27560
rect 2774 27548 2780 27560
rect 2832 27548 2838 27600
rect 7374 27548 7380 27600
rect 7432 27588 7438 27600
rect 7432 27560 8248 27588
rect 7432 27548 7438 27560
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 2866 27520 2872 27532
rect 1995 27492 2872 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 2866 27480 2872 27492
rect 2924 27480 2930 27532
rect 6632 27523 6690 27529
rect 6632 27489 6644 27523
rect 6678 27520 6690 27523
rect 7650 27520 7656 27532
rect 6678 27492 7656 27520
rect 6678 27489 6690 27492
rect 6632 27483 6690 27489
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 8220 27529 8248 27560
rect 9858 27548 9864 27600
rect 9916 27588 9922 27600
rect 10321 27591 10379 27597
rect 10321 27588 10333 27591
rect 9916 27560 10333 27588
rect 9916 27548 9922 27560
rect 10321 27557 10333 27560
rect 10367 27588 10379 27591
rect 10888 27588 10916 27628
rect 12250 27616 12256 27628
rect 12308 27616 12314 27668
rect 15102 27656 15108 27668
rect 14752 27628 15108 27656
rect 10367 27560 10916 27588
rect 10367 27557 10379 27560
rect 10321 27551 10379 27557
rect 10962 27548 10968 27600
rect 11020 27588 11026 27600
rect 14274 27588 14280 27600
rect 11020 27560 14280 27588
rect 11020 27548 11026 27560
rect 14274 27548 14280 27560
rect 14332 27548 14338 27600
rect 8205 27523 8263 27529
rect 8205 27489 8217 27523
rect 8251 27489 8263 27523
rect 8205 27483 8263 27489
rect 9493 27523 9551 27529
rect 9493 27489 9505 27523
rect 9539 27520 9551 27523
rect 9766 27520 9772 27532
rect 9539 27492 9772 27520
rect 9539 27489 9551 27492
rect 9493 27483 9551 27489
rect 9766 27480 9772 27492
rect 9824 27480 9830 27532
rect 10137 27523 10195 27529
rect 10137 27489 10149 27523
rect 10183 27489 10195 27523
rect 10137 27483 10195 27489
rect 10413 27523 10471 27529
rect 10413 27489 10425 27523
rect 10459 27489 10471 27523
rect 10413 27483 10471 27489
rect 5166 27412 5172 27464
rect 5224 27452 5230 27464
rect 6365 27455 6423 27461
rect 6365 27452 6377 27455
rect 5224 27424 6377 27452
rect 5224 27412 5230 27424
rect 6365 27421 6377 27424
rect 6411 27421 6423 27455
rect 6365 27415 6423 27421
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 10152 27452 10180 27483
rect 9456 27424 10180 27452
rect 10428 27452 10456 27483
rect 10502 27480 10508 27532
rect 10560 27520 10566 27532
rect 12152 27523 12210 27529
rect 10560 27492 10605 27520
rect 10560 27480 10566 27492
rect 12152 27489 12164 27523
rect 12198 27520 12210 27523
rect 12618 27520 12624 27532
rect 12198 27492 12624 27520
rect 12198 27489 12210 27492
rect 12152 27483 12210 27489
rect 12618 27480 12624 27492
rect 12676 27480 12682 27532
rect 13354 27480 13360 27532
rect 13412 27520 13418 27532
rect 14752 27529 14780 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 15286 27656 15292 27668
rect 15247 27628 15292 27656
rect 15286 27616 15292 27628
rect 15344 27616 15350 27668
rect 16022 27616 16028 27668
rect 16080 27656 16086 27668
rect 16301 27659 16359 27665
rect 16301 27656 16313 27659
rect 16080 27628 16313 27656
rect 16080 27616 16086 27628
rect 16301 27625 16313 27628
rect 16347 27625 16359 27659
rect 18046 27656 18052 27668
rect 18007 27628 18052 27656
rect 16301 27619 16359 27625
rect 18046 27616 18052 27628
rect 18104 27616 18110 27668
rect 15013 27591 15071 27597
rect 15013 27557 15025 27591
rect 15059 27588 15071 27591
rect 15378 27588 15384 27600
rect 15059 27560 15384 27588
rect 15059 27557 15071 27560
rect 15013 27551 15071 27557
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 15562 27548 15568 27600
rect 15620 27588 15626 27600
rect 15933 27591 15991 27597
rect 15933 27588 15945 27591
rect 15620 27560 15945 27588
rect 15620 27548 15626 27560
rect 15933 27557 15945 27560
rect 15979 27557 15991 27591
rect 16390 27588 16396 27600
rect 15933 27551 15991 27557
rect 16040 27560 16396 27588
rect 14737 27523 14795 27529
rect 14737 27520 14749 27523
rect 13412 27492 14749 27520
rect 13412 27480 13418 27492
rect 14737 27489 14749 27492
rect 14783 27489 14795 27523
rect 14737 27483 14795 27489
rect 14921 27523 14979 27529
rect 14921 27489 14933 27523
rect 14967 27489 14979 27523
rect 15102 27520 15108 27532
rect 15063 27492 15108 27520
rect 14921 27483 14979 27489
rect 11054 27452 11060 27464
rect 10428 27424 11060 27452
rect 9456 27412 9462 27424
rect 11054 27412 11060 27424
rect 11112 27412 11118 27464
rect 11882 27452 11888 27464
rect 11843 27424 11888 27452
rect 11882 27412 11888 27424
rect 11940 27412 11946 27464
rect 14366 27412 14372 27464
rect 14424 27452 14430 27464
rect 14936 27452 14964 27483
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 15194 27480 15200 27532
rect 15252 27520 15258 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 15252 27492 15761 27520
rect 15252 27480 15258 27492
rect 15749 27489 15761 27492
rect 15795 27520 15807 27523
rect 15838 27520 15844 27532
rect 15795 27492 15844 27520
rect 15795 27489 15807 27492
rect 15749 27483 15807 27489
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 16040 27529 16068 27560
rect 16390 27548 16396 27560
rect 16448 27548 16454 27600
rect 17402 27548 17408 27600
rect 17460 27588 17466 27600
rect 17681 27591 17739 27597
rect 17681 27588 17693 27591
rect 17460 27560 17693 27588
rect 17460 27548 17466 27560
rect 17681 27557 17693 27560
rect 17727 27557 17739 27591
rect 17681 27551 17739 27557
rect 17773 27591 17831 27597
rect 17773 27557 17785 27591
rect 17819 27588 17831 27591
rect 18322 27588 18328 27600
rect 17819 27560 18328 27588
rect 17819 27557 17831 27560
rect 17773 27551 17831 27557
rect 18322 27548 18328 27560
rect 18380 27588 18386 27600
rect 18874 27588 18880 27600
rect 18380 27560 18880 27588
rect 18380 27548 18386 27560
rect 18874 27548 18880 27560
rect 18932 27548 18938 27600
rect 20616 27591 20674 27597
rect 20616 27557 20628 27591
rect 20662 27588 20674 27591
rect 20806 27588 20812 27600
rect 20662 27560 20812 27588
rect 20662 27557 20674 27560
rect 20616 27551 20674 27557
rect 20806 27548 20812 27560
rect 20864 27548 20870 27600
rect 25774 27588 25780 27600
rect 25735 27560 25780 27588
rect 25774 27548 25780 27560
rect 25832 27548 25838 27600
rect 26050 27548 26056 27600
rect 26108 27588 26114 27600
rect 26513 27591 26571 27597
rect 26513 27588 26525 27591
rect 26108 27560 26525 27588
rect 26108 27548 26114 27560
rect 26513 27557 26525 27560
rect 26559 27557 26571 27591
rect 26513 27551 26571 27557
rect 16025 27523 16083 27529
rect 16025 27489 16037 27523
rect 16071 27489 16083 27523
rect 16025 27483 16083 27489
rect 16117 27523 16175 27529
rect 16117 27489 16129 27523
rect 16163 27489 16175 27523
rect 16117 27483 16175 27489
rect 15120 27452 15148 27480
rect 16132 27452 16160 27483
rect 16574 27480 16580 27532
rect 16632 27520 16638 27532
rect 16761 27523 16819 27529
rect 16761 27520 16773 27523
rect 16632 27492 16773 27520
rect 16632 27480 16638 27492
rect 16761 27489 16773 27492
rect 16807 27489 16819 27523
rect 16761 27483 16819 27489
rect 17497 27523 17555 27529
rect 17497 27489 17509 27523
rect 17543 27520 17555 27523
rect 17865 27523 17923 27529
rect 17543 27492 17724 27520
rect 17543 27489 17555 27492
rect 17497 27483 17555 27489
rect 17696 27464 17724 27492
rect 17865 27489 17877 27523
rect 17911 27520 17923 27523
rect 17954 27520 17960 27532
rect 17911 27492 17960 27520
rect 17911 27489 17923 27492
rect 17865 27483 17923 27489
rect 17954 27480 17960 27492
rect 18012 27480 18018 27532
rect 18414 27480 18420 27532
rect 18472 27520 18478 27532
rect 18509 27523 18567 27529
rect 18509 27520 18521 27523
rect 18472 27492 18521 27520
rect 18472 27480 18478 27492
rect 18509 27489 18521 27492
rect 18555 27489 18567 27523
rect 18509 27483 18567 27489
rect 24302 27480 24308 27532
rect 24360 27520 24366 27532
rect 25593 27523 25651 27529
rect 25593 27520 25605 27523
rect 24360 27492 25605 27520
rect 24360 27480 24366 27492
rect 25593 27489 25605 27492
rect 25639 27489 25651 27523
rect 25593 27483 25651 27489
rect 26329 27523 26387 27529
rect 26329 27489 26341 27523
rect 26375 27489 26387 27523
rect 26329 27483 26387 27489
rect 14424 27424 15056 27452
rect 15120 27424 16160 27452
rect 14424 27412 14430 27424
rect 7558 27344 7564 27396
rect 7616 27384 7622 27396
rect 15028 27384 15056 27424
rect 17678 27412 17684 27464
rect 17736 27412 17742 27464
rect 20346 27452 20352 27464
rect 20307 27424 20352 27452
rect 20346 27412 20352 27424
rect 20404 27412 20410 27464
rect 26344 27452 26372 27483
rect 26418 27480 26424 27532
rect 26476 27520 26482 27532
rect 26973 27523 27031 27529
rect 26973 27520 26985 27523
rect 26476 27492 26985 27520
rect 26476 27480 26482 27492
rect 26973 27489 26985 27492
rect 27019 27520 27031 27523
rect 27338 27520 27344 27532
rect 27019 27492 27344 27520
rect 27019 27489 27031 27492
rect 26973 27483 27031 27489
rect 27338 27480 27344 27492
rect 27396 27480 27402 27532
rect 26510 27452 26516 27464
rect 26344 27424 26516 27452
rect 26510 27412 26516 27424
rect 26568 27412 26574 27464
rect 17494 27384 17500 27396
rect 7616 27356 9720 27384
rect 15028 27356 17500 27384
rect 7616 27344 7622 27356
rect 1765 27319 1823 27325
rect 1765 27285 1777 27319
rect 1811 27316 1823 27319
rect 2958 27316 2964 27328
rect 1811 27288 2964 27316
rect 1811 27285 1823 27288
rect 1765 27279 1823 27285
rect 2958 27276 2964 27288
rect 3016 27276 3022 27328
rect 7374 27276 7380 27328
rect 7432 27316 7438 27328
rect 7745 27319 7803 27325
rect 7745 27316 7757 27319
rect 7432 27288 7757 27316
rect 7432 27276 7438 27288
rect 7745 27285 7757 27288
rect 7791 27285 7803 27319
rect 7745 27279 7803 27285
rect 8662 27276 8668 27328
rect 8720 27316 8726 27328
rect 9585 27319 9643 27325
rect 9585 27316 9597 27319
rect 8720 27288 9597 27316
rect 8720 27276 8726 27288
rect 9585 27285 9597 27288
rect 9631 27285 9643 27319
rect 9692 27316 9720 27356
rect 17494 27344 17500 27356
rect 17552 27344 17558 27396
rect 21726 27384 21732 27396
rect 21687 27356 21732 27384
rect 21726 27344 21732 27356
rect 21784 27344 21790 27396
rect 13078 27316 13084 27328
rect 9692 27288 13084 27316
rect 9585 27279 9643 27285
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 13262 27316 13268 27328
rect 13223 27288 13268 27316
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 16942 27316 16948 27328
rect 16903 27288 16948 27316
rect 16942 27276 16948 27288
rect 17000 27276 17006 27328
rect 18690 27316 18696 27328
rect 18651 27288 18696 27316
rect 18690 27276 18696 27288
rect 18748 27276 18754 27328
rect 1104 27226 28428 27248
rect 1104 27174 5536 27226
rect 5588 27174 5600 27226
rect 5652 27174 5664 27226
rect 5716 27174 5728 27226
rect 5780 27174 14644 27226
rect 14696 27174 14708 27226
rect 14760 27174 14772 27226
rect 14824 27174 14836 27226
rect 14888 27174 23752 27226
rect 23804 27174 23816 27226
rect 23868 27174 23880 27226
rect 23932 27174 23944 27226
rect 23996 27174 28428 27226
rect 1104 27152 28428 27174
rect 7650 27112 7656 27124
rect 7611 27084 7656 27112
rect 7650 27072 7656 27084
rect 7708 27072 7714 27124
rect 8665 27115 8723 27121
rect 8665 27081 8677 27115
rect 8711 27112 8723 27115
rect 8754 27112 8760 27124
rect 8711 27084 8760 27112
rect 8711 27081 8723 27084
rect 8665 27075 8723 27081
rect 8754 27072 8760 27084
rect 8812 27072 8818 27124
rect 9493 27115 9551 27121
rect 9493 27081 9505 27115
rect 9539 27112 9551 27115
rect 18690 27112 18696 27124
rect 9539 27084 18696 27112
rect 9539 27081 9551 27084
rect 9493 27075 9551 27081
rect 18690 27072 18696 27084
rect 18748 27072 18754 27124
rect 9858 27044 9864 27056
rect 9646 27016 9864 27044
rect 7116 26948 8156 26976
rect 7116 26920 7144 26948
rect 2130 26908 2136 26920
rect 2091 26880 2136 26908
rect 2130 26868 2136 26880
rect 2188 26868 2194 26920
rect 7098 26908 7104 26920
rect 7059 26880 7104 26908
rect 7098 26868 7104 26880
rect 7156 26868 7162 26920
rect 7374 26908 7380 26920
rect 7335 26880 7380 26908
rect 7374 26868 7380 26880
rect 7432 26868 7438 26920
rect 7469 26911 7527 26917
rect 7469 26877 7481 26911
rect 7515 26908 7527 26911
rect 7834 26908 7840 26920
rect 7515 26880 7840 26908
rect 7515 26877 7527 26880
rect 7469 26871 7527 26877
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 8128 26917 8156 26948
rect 9214 26936 9220 26988
rect 9272 26976 9278 26988
rect 9646 26976 9674 27016
rect 9858 27004 9864 27016
rect 9916 27004 9922 27056
rect 10042 27004 10048 27056
rect 10100 27044 10106 27056
rect 10597 27047 10655 27053
rect 10597 27044 10609 27047
rect 10100 27016 10609 27044
rect 10100 27004 10106 27016
rect 10597 27013 10609 27016
rect 10643 27013 10655 27047
rect 16390 27044 16396 27056
rect 10597 27007 10655 27013
rect 16132 27016 16396 27044
rect 15562 26976 15568 26988
rect 9272 26948 9674 26976
rect 9784 26948 12204 26976
rect 9272 26936 9278 26948
rect 8113 26911 8171 26917
rect 8113 26877 8125 26911
rect 8159 26877 8171 26911
rect 8481 26911 8539 26917
rect 8481 26908 8493 26911
rect 8113 26871 8171 26877
rect 8220 26880 8493 26908
rect 7285 26843 7343 26849
rect 7285 26809 7297 26843
rect 7331 26840 7343 26843
rect 7558 26840 7564 26852
rect 7331 26812 7564 26840
rect 7331 26809 7343 26812
rect 7285 26803 7343 26809
rect 7558 26800 7564 26812
rect 7616 26800 7622 26852
rect 7852 26840 7880 26868
rect 8220 26840 8248 26880
rect 8481 26877 8493 26880
rect 8527 26877 8539 26911
rect 8481 26871 8539 26877
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 9456 26880 9597 26908
rect 9456 26868 9462 26880
rect 9585 26877 9597 26880
rect 9631 26908 9643 26911
rect 9784 26908 9812 26948
rect 9631 26880 9812 26908
rect 9861 26911 9919 26917
rect 9631 26877 9643 26880
rect 9585 26871 9643 26877
rect 9861 26877 9873 26911
rect 9907 26877 9919 26911
rect 9861 26871 9919 26877
rect 9953 26911 10011 26917
rect 9953 26877 9965 26911
rect 9999 26877 10011 26911
rect 9953 26871 10011 26877
rect 7852 26812 8248 26840
rect 8297 26843 8355 26849
rect 8297 26809 8309 26843
rect 8343 26809 8355 26843
rect 8297 26803 8355 26809
rect 8389 26843 8447 26849
rect 8389 26809 8401 26843
rect 8435 26840 8447 26843
rect 9674 26840 9680 26852
rect 8435 26812 9680 26840
rect 8435 26809 8447 26812
rect 8389 26803 8447 26809
rect 8312 26772 8340 26803
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 9769 26843 9827 26849
rect 9769 26809 9781 26843
rect 9815 26809 9827 26843
rect 9769 26803 9827 26809
rect 9493 26775 9551 26781
rect 9493 26772 9505 26775
rect 8312 26744 9505 26772
rect 9493 26741 9505 26744
rect 9539 26741 9551 26775
rect 9493 26735 9551 26741
rect 9582 26732 9588 26784
rect 9640 26772 9646 26784
rect 9784 26772 9812 26803
rect 9867 26784 9895 26871
rect 9968 26840 9996 26871
rect 10134 26868 10140 26920
rect 10192 26908 10198 26920
rect 10781 26911 10839 26917
rect 10781 26908 10793 26911
rect 10192 26880 10793 26908
rect 10192 26868 10198 26880
rect 10781 26877 10793 26880
rect 10827 26877 10839 26911
rect 10781 26871 10839 26877
rect 11882 26868 11888 26920
rect 11940 26908 11946 26920
rect 12069 26911 12127 26917
rect 12069 26908 12081 26911
rect 11940 26880 12081 26908
rect 11940 26868 11946 26880
rect 12069 26877 12081 26880
rect 12115 26877 12127 26911
rect 12176 26908 12204 26948
rect 15212 26948 15568 26976
rect 13354 26908 13360 26920
rect 12176 26880 13360 26908
rect 12069 26871 12127 26877
rect 13354 26868 13360 26880
rect 13412 26868 13418 26920
rect 13909 26911 13967 26917
rect 13909 26908 13921 26911
rect 13464 26880 13921 26908
rect 10502 26840 10508 26852
rect 9968 26812 10508 26840
rect 10502 26800 10508 26812
rect 10560 26800 10566 26852
rect 12336 26843 12394 26849
rect 12336 26809 12348 26843
rect 12382 26840 12394 26843
rect 12710 26840 12716 26852
rect 12382 26812 12716 26840
rect 12382 26809 12394 26812
rect 12336 26803 12394 26809
rect 12710 26800 12716 26812
rect 12768 26800 12774 26852
rect 9640 26744 9812 26772
rect 9640 26732 9646 26744
rect 9854 26732 9860 26784
rect 9912 26732 9918 26784
rect 9950 26732 9956 26784
rect 10008 26772 10014 26784
rect 10137 26775 10195 26781
rect 10137 26772 10149 26775
rect 10008 26744 10149 26772
rect 10008 26732 10014 26744
rect 10137 26741 10149 26744
rect 10183 26741 10195 26775
rect 10137 26735 10195 26741
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 13464 26781 13492 26880
rect 13909 26877 13921 26880
rect 13955 26877 13967 26911
rect 13909 26871 13967 26877
rect 15013 26911 15071 26917
rect 15013 26877 15025 26911
rect 15059 26908 15071 26911
rect 15102 26908 15108 26920
rect 15059 26880 15108 26908
rect 15059 26877 15071 26880
rect 15013 26871 15071 26877
rect 15102 26868 15108 26880
rect 15160 26868 15166 26920
rect 15212 26917 15240 26948
rect 15562 26936 15568 26948
rect 15620 26976 15626 26988
rect 16022 26976 16028 26988
rect 15620 26948 16028 26976
rect 15620 26936 15626 26948
rect 16022 26936 16028 26948
rect 16080 26936 16086 26988
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26877 15255 26911
rect 15197 26871 15255 26877
rect 15381 26911 15439 26917
rect 15381 26877 15393 26911
rect 15427 26908 15439 26911
rect 15470 26908 15476 26920
rect 15427 26880 15476 26908
rect 15427 26877 15439 26880
rect 15381 26871 15439 26877
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 16132 26917 16160 27016
rect 16390 27004 16396 27016
rect 16448 27004 16454 27056
rect 26878 27044 26884 27056
rect 26839 27016 26884 27044
rect 26878 27004 26884 27016
rect 26936 27004 26942 27056
rect 16206 26936 16212 26988
rect 16264 26976 16270 26988
rect 16264 26948 17724 26976
rect 16264 26936 16270 26948
rect 16117 26911 16175 26917
rect 16117 26877 16129 26911
rect 16163 26877 16175 26911
rect 16117 26871 16175 26877
rect 16390 26868 16396 26920
rect 16448 26908 16454 26920
rect 17313 26911 17371 26917
rect 17313 26908 17325 26911
rect 16448 26880 17325 26908
rect 16448 26868 16454 26880
rect 17313 26877 17325 26880
rect 17359 26877 17371 26911
rect 17494 26908 17500 26920
rect 17455 26880 17500 26908
rect 17313 26871 17371 26877
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 17696 26917 17724 26948
rect 17681 26911 17739 26917
rect 17681 26877 17693 26911
rect 17727 26877 17739 26911
rect 18322 26908 18328 26920
rect 18283 26880 18328 26908
rect 17681 26871 17739 26877
rect 18322 26868 18328 26880
rect 18380 26868 18386 26920
rect 18782 26868 18788 26920
rect 18840 26908 18846 26920
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 18840 26880 18981 26908
rect 18840 26868 18846 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 18969 26871 19027 26877
rect 21453 26911 21511 26917
rect 21453 26877 21465 26911
rect 21499 26908 21511 26911
rect 21726 26908 21732 26920
rect 21499 26880 21732 26908
rect 21499 26877 21511 26880
rect 21453 26871 21511 26877
rect 21726 26868 21732 26880
rect 21784 26868 21790 26920
rect 21818 26868 21824 26920
rect 21876 26908 21882 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 21876 26880 22845 26908
rect 21876 26868 21882 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 22833 26871 22891 26877
rect 22922 26868 22928 26920
rect 22980 26908 22986 26920
rect 23109 26911 23167 26917
rect 23109 26908 23121 26911
rect 22980 26880 23121 26908
rect 22980 26868 22986 26880
rect 23109 26877 23121 26880
rect 23155 26877 23167 26911
rect 23109 26871 23167 26877
rect 23201 26911 23259 26917
rect 23201 26877 23213 26911
rect 23247 26908 23259 26911
rect 24302 26908 24308 26920
rect 23247 26880 24308 26908
rect 23247 26877 23259 26880
rect 23201 26871 23259 26877
rect 24302 26868 24308 26880
rect 24360 26868 24366 26920
rect 15289 26843 15347 26849
rect 15289 26809 15301 26843
rect 15335 26840 15347 26843
rect 16666 26840 16672 26852
rect 15335 26812 16672 26840
rect 15335 26809 15347 26812
rect 15289 26803 15347 26809
rect 16666 26800 16672 26812
rect 16724 26800 16730 26852
rect 17589 26843 17647 26849
rect 17589 26809 17601 26843
rect 17635 26840 17647 26843
rect 18230 26840 18236 26852
rect 17635 26812 18236 26840
rect 17635 26809 17647 26812
rect 17589 26803 17647 26809
rect 18230 26800 18236 26812
rect 18288 26800 18294 26852
rect 23017 26843 23075 26849
rect 23017 26809 23029 26843
rect 23063 26809 23075 26843
rect 23017 26803 23075 26809
rect 13449 26775 13507 26781
rect 13449 26772 13461 26775
rect 12584 26744 13461 26772
rect 12584 26732 12590 26744
rect 13449 26741 13461 26744
rect 13495 26741 13507 26775
rect 13449 26735 13507 26741
rect 14001 26775 14059 26781
rect 14001 26741 14013 26775
rect 14047 26772 14059 26775
rect 14182 26772 14188 26784
rect 14047 26744 14188 26772
rect 14047 26741 14059 26744
rect 14001 26735 14059 26741
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 15562 26772 15568 26784
rect 15523 26744 15568 26772
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 16209 26775 16267 26781
rect 16209 26741 16221 26775
rect 16255 26772 16267 26775
rect 16574 26772 16580 26784
rect 16255 26744 16580 26772
rect 16255 26741 16267 26744
rect 16209 26735 16267 26741
rect 16574 26732 16580 26744
rect 16632 26732 16638 26784
rect 17862 26772 17868 26784
rect 17823 26744 17868 26772
rect 17862 26732 17868 26744
rect 17920 26732 17926 26784
rect 18417 26775 18475 26781
rect 18417 26741 18429 26775
rect 18463 26772 18475 26775
rect 18506 26772 18512 26784
rect 18463 26744 18512 26772
rect 18463 26741 18475 26744
rect 18417 26735 18475 26741
rect 18506 26732 18512 26744
rect 18564 26732 18570 26784
rect 18598 26732 18604 26784
rect 18656 26772 18662 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 18656 26744 19073 26772
rect 18656 26732 18662 26744
rect 19061 26741 19073 26744
rect 19107 26741 19119 26775
rect 21542 26772 21548 26784
rect 21503 26744 21548 26772
rect 19061 26735 19119 26741
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 23032 26772 23060 26803
rect 23290 26800 23296 26852
rect 23348 26840 23354 26852
rect 26697 26843 26755 26849
rect 26697 26840 26709 26843
rect 23348 26812 26709 26840
rect 23348 26800 23354 26812
rect 26697 26809 26709 26812
rect 26743 26809 26755 26843
rect 26697 26803 26755 26809
rect 23198 26772 23204 26784
rect 23032 26744 23204 26772
rect 23198 26732 23204 26744
rect 23256 26732 23262 26784
rect 23382 26772 23388 26784
rect 23343 26744 23388 26772
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 1104 26682 28428 26704
rect 1104 26630 10090 26682
rect 10142 26630 10154 26682
rect 10206 26630 10218 26682
rect 10270 26630 10282 26682
rect 10334 26630 19198 26682
rect 19250 26630 19262 26682
rect 19314 26630 19326 26682
rect 19378 26630 19390 26682
rect 19442 26630 28428 26682
rect 1104 26608 28428 26630
rect 1946 26568 1952 26580
rect 1907 26540 1952 26568
rect 1946 26528 1952 26540
rect 2004 26528 2010 26580
rect 9490 26528 9496 26580
rect 9548 26568 9554 26580
rect 16485 26571 16543 26577
rect 9548 26540 10456 26568
rect 9548 26528 9554 26540
rect 9760 26503 9818 26509
rect 9760 26469 9772 26503
rect 9806 26500 9818 26503
rect 9950 26500 9956 26512
rect 9806 26472 9956 26500
rect 9806 26469 9818 26472
rect 9760 26463 9818 26469
rect 9950 26460 9956 26472
rect 10008 26460 10014 26512
rect 10428 26500 10456 26540
rect 16485 26537 16497 26571
rect 16531 26568 16543 26571
rect 16666 26568 16672 26580
rect 16531 26540 16672 26568
rect 16531 26537 16543 26540
rect 16485 26531 16543 26537
rect 16666 26528 16672 26540
rect 16724 26528 16730 26580
rect 18230 26528 18236 26580
rect 18288 26568 18294 26580
rect 18509 26571 18567 26577
rect 18509 26568 18521 26571
rect 18288 26540 18521 26568
rect 18288 26528 18294 26540
rect 18509 26537 18521 26540
rect 18555 26568 18567 26571
rect 18782 26568 18788 26580
rect 18555 26540 18788 26568
rect 18555 26537 18567 26540
rect 18509 26531 18567 26537
rect 18782 26528 18788 26540
rect 18840 26528 18846 26580
rect 22278 26568 22284 26580
rect 22191 26540 22284 26568
rect 22278 26528 22284 26540
rect 22336 26568 22342 26580
rect 23290 26568 23296 26580
rect 22336 26540 23296 26568
rect 22336 26528 22342 26540
rect 23290 26528 23296 26540
rect 23348 26528 23354 26580
rect 24302 26568 24308 26580
rect 24263 26540 24308 26568
rect 24302 26528 24308 26540
rect 24360 26528 24366 26580
rect 11882 26500 11888 26512
rect 10428 26472 11888 26500
rect 1857 26435 1915 26441
rect 1857 26401 1869 26435
rect 1903 26432 1915 26435
rect 2130 26432 2136 26444
rect 1903 26404 2136 26432
rect 1903 26401 1915 26404
rect 1857 26395 1915 26401
rect 2130 26392 2136 26404
rect 2188 26432 2194 26444
rect 11054 26432 11060 26444
rect 2188 26404 11060 26432
rect 2188 26392 2194 26404
rect 11054 26392 11060 26404
rect 11112 26392 11118 26444
rect 11808 26441 11836 26472
rect 11882 26460 11888 26472
rect 11940 26460 11946 26512
rect 12060 26503 12118 26509
rect 12060 26469 12072 26503
rect 12106 26500 12118 26503
rect 13722 26500 13728 26512
rect 12106 26472 13728 26500
rect 12106 26469 12118 26472
rect 12060 26463 12118 26469
rect 13722 26460 13728 26472
rect 13780 26460 13786 26512
rect 15372 26503 15430 26509
rect 15372 26469 15384 26503
rect 15418 26500 15430 26503
rect 15562 26500 15568 26512
rect 15418 26472 15568 26500
rect 15418 26469 15430 26472
rect 15372 26463 15430 26469
rect 15562 26460 15568 26472
rect 15620 26460 15626 26512
rect 17396 26503 17454 26509
rect 17396 26469 17408 26503
rect 17442 26500 17454 26503
rect 17862 26500 17868 26512
rect 17442 26472 17868 26500
rect 17442 26469 17454 26472
rect 17396 26463 17454 26469
rect 17862 26460 17868 26472
rect 17920 26460 17926 26512
rect 23192 26503 23250 26509
rect 23192 26469 23204 26503
rect 23238 26500 23250 26503
rect 23382 26500 23388 26512
rect 23238 26472 23388 26500
rect 23238 26469 23250 26472
rect 23192 26463 23250 26469
rect 23382 26460 23388 26472
rect 23440 26460 23446 26512
rect 26789 26503 26847 26509
rect 26789 26469 26801 26503
rect 26835 26500 26847 26503
rect 27430 26500 27436 26512
rect 26835 26472 27436 26500
rect 26835 26469 26847 26472
rect 26789 26463 26847 26469
rect 27430 26460 27436 26472
rect 27488 26460 27494 26512
rect 27706 26500 27712 26512
rect 27667 26472 27712 26500
rect 27706 26460 27712 26472
rect 27764 26460 27770 26512
rect 11793 26435 11851 26441
rect 11793 26401 11805 26435
rect 11839 26401 11851 26435
rect 13262 26432 13268 26444
rect 11793 26395 11851 26401
rect 13004 26404 13268 26432
rect 9490 26364 9496 26376
rect 9451 26336 9496 26364
rect 9490 26324 9496 26336
rect 9548 26324 9554 26376
rect 2130 26188 2136 26240
rect 2188 26228 2194 26240
rect 9858 26228 9864 26240
rect 2188 26200 9864 26228
rect 2188 26188 2194 26200
rect 9858 26188 9864 26200
rect 9916 26228 9922 26240
rect 10873 26231 10931 26237
rect 10873 26228 10885 26231
rect 9916 26200 10885 26228
rect 9916 26188 9922 26200
rect 10873 26197 10885 26200
rect 10919 26197 10931 26231
rect 10873 26191 10931 26197
rect 12158 26188 12164 26240
rect 12216 26228 12222 26240
rect 13004 26228 13032 26404
rect 13262 26392 13268 26404
rect 13320 26432 13326 26444
rect 13633 26435 13691 26441
rect 13633 26432 13645 26435
rect 13320 26404 13645 26432
rect 13320 26392 13326 26404
rect 13633 26401 13645 26404
rect 13679 26401 13691 26435
rect 13633 26395 13691 26401
rect 14458 26392 14464 26444
rect 14516 26432 14522 26444
rect 15105 26435 15163 26441
rect 15105 26432 15117 26435
rect 14516 26404 15117 26432
rect 14516 26392 14522 26404
rect 15105 26401 15117 26404
rect 15151 26432 15163 26435
rect 17129 26435 17187 26441
rect 17129 26432 17141 26435
rect 15151 26404 17141 26432
rect 15151 26401 15163 26404
rect 15105 26395 15163 26401
rect 17129 26401 17141 26404
rect 17175 26432 17187 26435
rect 17218 26432 17224 26444
rect 17175 26404 17224 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 17218 26392 17224 26404
rect 17276 26432 17282 26444
rect 20346 26432 20352 26444
rect 17276 26404 20352 26432
rect 17276 26392 17282 26404
rect 20346 26392 20352 26404
rect 20404 26432 20410 26444
rect 20901 26435 20959 26441
rect 20901 26432 20913 26435
rect 20404 26404 20913 26432
rect 20404 26392 20410 26404
rect 20901 26401 20913 26404
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 21168 26435 21226 26441
rect 21168 26401 21180 26435
rect 21214 26432 21226 26435
rect 21450 26432 21456 26444
rect 21214 26404 21456 26432
rect 21214 26401 21226 26404
rect 21168 26395 21226 26401
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 27154 26392 27160 26444
rect 27212 26432 27218 26444
rect 27525 26435 27583 26441
rect 27525 26432 27537 26435
rect 27212 26404 27537 26432
rect 27212 26392 27218 26404
rect 27525 26401 27537 26404
rect 27571 26401 27583 26435
rect 27525 26395 27583 26401
rect 22830 26324 22836 26376
rect 22888 26364 22894 26376
rect 22925 26367 22983 26373
rect 22925 26364 22937 26367
rect 22888 26336 22937 26364
rect 22888 26324 22894 26336
rect 22925 26333 22937 26336
rect 22971 26333 22983 26367
rect 22925 26327 22983 26333
rect 13725 26299 13783 26305
rect 13725 26265 13737 26299
rect 13771 26296 13783 26299
rect 14458 26296 14464 26308
rect 13771 26268 14464 26296
rect 13771 26265 13783 26268
rect 13725 26259 13783 26265
rect 14458 26256 14464 26268
rect 14516 26256 14522 26308
rect 26970 26296 26976 26308
rect 26931 26268 26976 26296
rect 26970 26256 26976 26268
rect 27028 26256 27034 26308
rect 13170 26228 13176 26240
rect 12216 26200 13032 26228
rect 13131 26200 13176 26228
rect 12216 26188 12222 26200
rect 13170 26188 13176 26200
rect 13228 26188 13234 26240
rect 1104 26138 28428 26160
rect 1104 26086 5536 26138
rect 5588 26086 5600 26138
rect 5652 26086 5664 26138
rect 5716 26086 5728 26138
rect 5780 26086 14644 26138
rect 14696 26086 14708 26138
rect 14760 26086 14772 26138
rect 14824 26086 14836 26138
rect 14888 26086 23752 26138
rect 23804 26086 23816 26138
rect 23868 26086 23880 26138
rect 23932 26086 23944 26138
rect 23996 26086 28428 26138
rect 1104 26064 28428 26086
rect 7101 26027 7159 26033
rect 7101 25993 7113 26027
rect 7147 25993 7159 26027
rect 7101 25987 7159 25993
rect 7837 26027 7895 26033
rect 7837 25993 7849 26027
rect 7883 26024 7895 26027
rect 12342 26024 12348 26036
rect 7883 25996 12348 26024
rect 7883 25993 7895 25996
rect 7837 25987 7895 25993
rect 7116 25956 7144 25987
rect 12342 25984 12348 25996
rect 12400 25984 12406 26036
rect 12618 26024 12624 26036
rect 12579 25996 12624 26024
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 21450 26024 21456 26036
rect 14752 25996 18368 26024
rect 21411 25996 21456 26024
rect 8202 25956 8208 25968
rect 7116 25928 8208 25956
rect 8202 25916 8208 25928
rect 8260 25916 8266 25968
rect 14274 25916 14280 25968
rect 14332 25956 14338 25968
rect 14752 25965 14780 25996
rect 14737 25959 14795 25965
rect 14332 25928 14596 25956
rect 14332 25916 14338 25928
rect 1670 25888 1676 25900
rect 1631 25860 1676 25888
rect 1670 25848 1676 25860
rect 1728 25848 1734 25900
rect 5460 25860 9904 25888
rect 1489 25823 1547 25829
rect 1489 25789 1501 25823
rect 1535 25820 1547 25823
rect 2130 25820 2136 25832
rect 1535 25792 2136 25820
rect 1535 25789 1547 25792
rect 1489 25783 1547 25789
rect 2130 25780 2136 25792
rect 2188 25780 2194 25832
rect 2866 25820 2872 25832
rect 2827 25792 2872 25820
rect 2866 25780 2872 25792
rect 2924 25780 2930 25832
rect 5258 25820 5264 25832
rect 5219 25792 5264 25820
rect 5258 25780 5264 25792
rect 5316 25780 5322 25832
rect 5460 25829 5488 25860
rect 5445 25823 5503 25829
rect 5445 25789 5457 25823
rect 5491 25789 5503 25823
rect 5445 25783 5503 25789
rect 5629 25823 5687 25829
rect 5629 25789 5641 25823
rect 5675 25820 5687 25823
rect 5902 25820 5908 25832
rect 5675 25792 5908 25820
rect 5675 25789 5687 25792
rect 5629 25783 5687 25789
rect 5902 25780 5908 25792
rect 5960 25780 5966 25832
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25820 6883 25823
rect 7374 25820 7380 25832
rect 6871 25792 7380 25820
rect 6871 25789 6883 25792
rect 6825 25783 6883 25789
rect 7374 25780 7380 25792
rect 7432 25780 7438 25832
rect 7466 25780 7472 25832
rect 7524 25820 7530 25832
rect 7745 25823 7803 25829
rect 7745 25820 7757 25823
rect 7524 25792 7757 25820
rect 7524 25780 7530 25792
rect 7745 25789 7757 25792
rect 7791 25789 7803 25823
rect 7745 25783 7803 25789
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 9769 25823 9827 25829
rect 9769 25820 9781 25823
rect 9548 25792 9781 25820
rect 9548 25780 9554 25792
rect 9769 25789 9781 25792
rect 9815 25789 9827 25823
rect 9876 25820 9904 25860
rect 11238 25848 11244 25900
rect 11296 25888 11302 25900
rect 14458 25888 14464 25900
rect 11296 25860 14320 25888
rect 14419 25860 14464 25888
rect 11296 25848 11302 25860
rect 10410 25820 10416 25832
rect 9876 25792 10416 25820
rect 9769 25783 9827 25789
rect 10410 25780 10416 25792
rect 10468 25780 10474 25832
rect 12066 25820 12072 25832
rect 12027 25792 12072 25820
rect 12066 25780 12072 25792
rect 12124 25780 12130 25832
rect 12158 25780 12164 25832
rect 12216 25820 12222 25832
rect 12452 25829 12480 25860
rect 12345 25823 12403 25829
rect 12345 25820 12357 25823
rect 12216 25792 12357 25820
rect 12216 25780 12222 25792
rect 12345 25789 12357 25792
rect 12391 25789 12403 25823
rect 12345 25783 12403 25789
rect 12437 25823 12495 25829
rect 12437 25789 12449 25823
rect 12483 25789 12495 25823
rect 12437 25783 12495 25789
rect 13541 25823 13599 25829
rect 13541 25789 13553 25823
rect 13587 25789 13599 25823
rect 13541 25783 13599 25789
rect 3136 25755 3194 25761
rect 3136 25721 3148 25755
rect 3182 25752 3194 25755
rect 3326 25752 3332 25764
rect 3182 25724 3332 25752
rect 3182 25721 3194 25724
rect 3136 25715 3194 25721
rect 3326 25712 3332 25724
rect 3384 25712 3390 25764
rect 5537 25755 5595 25761
rect 5537 25721 5549 25755
rect 5583 25752 5595 25755
rect 7484 25752 7512 25780
rect 5583 25724 7512 25752
rect 10036 25755 10094 25761
rect 5583 25721 5595 25724
rect 5537 25715 5595 25721
rect 10036 25721 10048 25755
rect 10082 25752 10094 25755
rect 11422 25752 11428 25764
rect 10082 25724 11428 25752
rect 10082 25721 10094 25724
rect 10036 25715 10094 25721
rect 11422 25712 11428 25724
rect 11480 25712 11486 25764
rect 12250 25712 12256 25764
rect 12308 25752 12314 25764
rect 13556 25752 13584 25783
rect 13630 25780 13636 25832
rect 13688 25820 13694 25832
rect 13817 25823 13875 25829
rect 13817 25820 13829 25823
rect 13688 25792 13829 25820
rect 13688 25780 13694 25792
rect 13817 25789 13829 25792
rect 13863 25789 13875 25823
rect 13817 25783 13875 25789
rect 14090 25780 14096 25832
rect 14148 25820 14154 25832
rect 14185 25823 14243 25829
rect 14185 25820 14197 25823
rect 14148 25792 14197 25820
rect 14148 25780 14154 25792
rect 14185 25789 14197 25792
rect 14231 25789 14243 25823
rect 14185 25783 14243 25789
rect 13998 25752 14004 25764
rect 12308 25724 12353 25752
rect 13556 25724 14004 25752
rect 12308 25712 12314 25724
rect 13998 25712 14004 25724
rect 14056 25712 14062 25764
rect 14292 25752 14320 25860
rect 14458 25848 14464 25860
rect 14516 25848 14522 25900
rect 14568 25888 14596 25928
rect 14737 25925 14749 25959
rect 14783 25925 14795 25959
rect 16390 25956 16396 25968
rect 14737 25919 14795 25925
rect 15856 25928 16396 25956
rect 15856 25888 15884 25928
rect 16390 25916 16396 25928
rect 16448 25916 16454 25968
rect 18340 25888 18368 25996
rect 21450 25984 21456 25996
rect 21508 25984 21514 26036
rect 24210 26024 24216 26036
rect 24171 25996 24216 26024
rect 24210 25984 24216 25996
rect 24268 25984 24274 26036
rect 26878 25888 26884 25900
rect 14568 25860 15884 25888
rect 14737 25823 14795 25829
rect 14737 25789 14749 25823
rect 14783 25820 14795 25823
rect 15654 25820 15660 25832
rect 14783 25792 15660 25820
rect 14783 25789 14795 25792
rect 14737 25783 14795 25789
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 15856 25829 15884 25860
rect 16132 25860 17448 25888
rect 18340 25860 22968 25888
rect 26839 25860 26884 25888
rect 15841 25823 15899 25829
rect 15841 25789 15853 25823
rect 15887 25789 15899 25823
rect 16022 25820 16028 25832
rect 15983 25792 16028 25820
rect 15841 25783 15899 25789
rect 16022 25780 16028 25792
rect 16080 25780 16086 25832
rect 16132 25829 16160 25860
rect 16117 25823 16175 25829
rect 16117 25789 16129 25823
rect 16163 25789 16175 25823
rect 16117 25783 16175 25789
rect 16206 25780 16212 25832
rect 16264 25820 16270 25832
rect 16264 25792 16309 25820
rect 16264 25780 16270 25792
rect 17218 25780 17224 25832
rect 17276 25820 17282 25832
rect 17313 25823 17371 25829
rect 17313 25820 17325 25823
rect 17276 25792 17325 25820
rect 17276 25780 17282 25792
rect 17313 25789 17325 25792
rect 17359 25789 17371 25823
rect 17420 25820 17448 25860
rect 20898 25820 20904 25832
rect 17420 25792 17908 25820
rect 20859 25792 20904 25820
rect 17313 25783 17371 25789
rect 16224 25752 16252 25780
rect 17558 25755 17616 25761
rect 17558 25752 17570 25755
rect 14292 25724 16252 25752
rect 16408 25724 17570 25752
rect 16040 25696 16068 25724
rect 4246 25684 4252 25696
rect 4207 25656 4252 25684
rect 4246 25644 4252 25656
rect 4304 25644 4310 25696
rect 5810 25684 5816 25696
rect 5771 25656 5816 25684
rect 5810 25644 5816 25656
rect 5868 25644 5874 25696
rect 6086 25644 6092 25696
rect 6144 25684 6150 25696
rect 7285 25687 7343 25693
rect 7285 25684 7297 25687
rect 6144 25656 7297 25684
rect 6144 25644 6150 25656
rect 7285 25653 7297 25656
rect 7331 25653 7343 25687
rect 11146 25684 11152 25696
rect 11107 25656 11152 25684
rect 7285 25647 7343 25653
rect 11146 25644 11152 25656
rect 11204 25644 11210 25696
rect 12618 25644 12624 25696
rect 12676 25684 12682 25696
rect 14274 25684 14280 25696
rect 12676 25656 14280 25684
rect 12676 25644 12682 25656
rect 14274 25644 14280 25656
rect 14332 25644 14338 25696
rect 16022 25644 16028 25696
rect 16080 25644 16086 25696
rect 16408 25693 16436 25724
rect 17558 25721 17570 25724
rect 17604 25721 17616 25755
rect 17558 25715 17616 25721
rect 16393 25687 16451 25693
rect 16393 25653 16405 25687
rect 16439 25653 16451 25687
rect 17880 25684 17908 25792
rect 20898 25780 20904 25792
rect 20956 25780 20962 25832
rect 21269 25823 21327 25829
rect 21269 25789 21281 25823
rect 21315 25820 21327 25823
rect 22278 25820 22284 25832
rect 21315 25792 22284 25820
rect 21315 25789 21327 25792
rect 21269 25783 21327 25789
rect 22278 25780 22284 25792
rect 22336 25780 22342 25832
rect 22830 25820 22836 25832
rect 22743 25792 22836 25820
rect 22830 25780 22836 25792
rect 22888 25780 22894 25832
rect 22940 25820 22968 25860
rect 26878 25848 26884 25860
rect 26936 25848 26942 25900
rect 24673 25823 24731 25829
rect 24673 25820 24685 25823
rect 22940 25792 24685 25820
rect 24673 25789 24685 25792
rect 24719 25789 24731 25823
rect 24673 25783 24731 25789
rect 25041 25823 25099 25829
rect 25041 25789 25053 25823
rect 25087 25820 25099 25823
rect 26602 25820 26608 25832
rect 25087 25792 26608 25820
rect 25087 25789 25099 25792
rect 25041 25783 25099 25789
rect 26602 25780 26608 25792
rect 26660 25820 26666 25832
rect 26697 25823 26755 25829
rect 26697 25820 26709 25823
rect 26660 25792 26709 25820
rect 26660 25780 26666 25792
rect 26697 25789 26709 25792
rect 26743 25789 26755 25823
rect 26697 25783 26755 25789
rect 21082 25752 21088 25764
rect 21043 25724 21088 25752
rect 21082 25712 21088 25724
rect 21140 25712 21146 25764
rect 21177 25755 21235 25761
rect 21177 25721 21189 25755
rect 21223 25752 21235 25755
rect 22848 25752 22876 25780
rect 23100 25755 23158 25761
rect 21223 25724 22094 25752
rect 22848 25724 23060 25752
rect 21223 25721 21235 25724
rect 21177 25715 21235 25721
rect 18693 25687 18751 25693
rect 18693 25684 18705 25687
rect 17880 25656 18705 25684
rect 16393 25647 16451 25653
rect 18693 25653 18705 25656
rect 18739 25684 18751 25687
rect 18874 25684 18880 25696
rect 18739 25656 18880 25684
rect 18739 25653 18751 25656
rect 18693 25647 18751 25653
rect 18874 25644 18880 25656
rect 18932 25644 18938 25696
rect 22066 25684 22094 25724
rect 22278 25684 22284 25696
rect 22066 25656 22284 25684
rect 22278 25644 22284 25656
rect 22336 25684 22342 25696
rect 22922 25684 22928 25696
rect 22336 25656 22928 25684
rect 22336 25644 22342 25656
rect 22922 25644 22928 25656
rect 22980 25644 22986 25696
rect 23032 25684 23060 25724
rect 23100 25721 23112 25755
rect 23146 25752 23158 25755
rect 23382 25752 23388 25764
rect 23146 25724 23388 25752
rect 23146 25721 23158 25724
rect 23100 25715 23158 25721
rect 23382 25712 23388 25724
rect 23440 25712 23446 25764
rect 24762 25712 24768 25764
rect 24820 25752 24826 25764
rect 24857 25755 24915 25761
rect 24857 25752 24869 25755
rect 24820 25724 24869 25752
rect 24820 25712 24826 25724
rect 24857 25721 24869 25724
rect 24903 25721 24915 25755
rect 24857 25715 24915 25721
rect 24946 25712 24952 25764
rect 25004 25752 25010 25764
rect 25004 25724 25049 25752
rect 25004 25712 25010 25724
rect 24118 25684 24124 25696
rect 23032 25656 24124 25684
rect 24118 25644 24124 25656
rect 24176 25644 24182 25696
rect 25222 25684 25228 25696
rect 25183 25656 25228 25684
rect 25222 25644 25228 25656
rect 25280 25644 25286 25696
rect 1104 25594 28428 25616
rect 1104 25542 10090 25594
rect 10142 25542 10154 25594
rect 10206 25542 10218 25594
rect 10270 25542 10282 25594
rect 10334 25542 19198 25594
rect 19250 25542 19262 25594
rect 19314 25542 19326 25594
rect 19378 25542 19390 25594
rect 19442 25542 28428 25594
rect 1104 25520 28428 25542
rect 3326 25480 3332 25492
rect 3287 25452 3332 25480
rect 3326 25440 3332 25452
rect 3384 25440 3390 25492
rect 4246 25440 4252 25492
rect 4304 25480 4310 25492
rect 6549 25483 6607 25489
rect 4304 25452 5939 25480
rect 4304 25440 4310 25452
rect 2958 25412 2964 25424
rect 2919 25384 2964 25412
rect 2958 25372 2964 25384
rect 3016 25372 3022 25424
rect 3053 25415 3111 25421
rect 3053 25381 3065 25415
rect 3099 25412 3111 25415
rect 4264 25412 4292 25440
rect 3099 25384 4292 25412
rect 5436 25415 5494 25421
rect 3099 25381 3111 25384
rect 3053 25375 3111 25381
rect 5436 25381 5448 25415
rect 5482 25412 5494 25415
rect 5810 25412 5816 25424
rect 5482 25384 5816 25412
rect 5482 25381 5494 25384
rect 5436 25375 5494 25381
rect 5810 25372 5816 25384
rect 5868 25372 5874 25424
rect 5911 25412 5939 25452
rect 6549 25449 6561 25483
rect 6595 25480 6607 25483
rect 7466 25480 7472 25492
rect 6595 25452 7472 25480
rect 6595 25449 6607 25452
rect 6549 25443 6607 25449
rect 7466 25440 7472 25452
rect 7524 25440 7530 25492
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 10870 25480 10876 25492
rect 9732 25452 10876 25480
rect 9732 25440 9738 25452
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 11422 25480 11428 25492
rect 11383 25452 11428 25480
rect 11422 25440 11428 25452
rect 11480 25440 11486 25492
rect 12250 25440 12256 25492
rect 12308 25440 12314 25492
rect 12710 25440 12716 25492
rect 12768 25480 12774 25492
rect 12805 25483 12863 25489
rect 12805 25480 12817 25483
rect 12768 25452 12817 25480
rect 12768 25440 12774 25452
rect 12805 25449 12817 25452
rect 12851 25449 12863 25483
rect 12805 25443 12863 25449
rect 13078 25440 13084 25492
rect 13136 25480 13142 25492
rect 13136 25452 13676 25480
rect 13136 25440 13142 25452
rect 11146 25412 11152 25424
rect 5911 25384 8156 25412
rect 1394 25344 1400 25356
rect 1355 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25304 1458 25356
rect 2777 25347 2835 25353
rect 2777 25313 2789 25347
rect 2823 25344 2835 25347
rect 3142 25344 3148 25356
rect 2823 25316 2857 25344
rect 3103 25316 3148 25344
rect 2823 25313 2835 25316
rect 2777 25307 2835 25313
rect 2682 25236 2688 25288
rect 2740 25276 2746 25288
rect 2792 25276 2820 25307
rect 3142 25304 3148 25316
rect 3200 25304 3206 25356
rect 3326 25304 3332 25356
rect 3384 25344 3390 25356
rect 4249 25347 4307 25353
rect 4249 25344 4261 25347
rect 3384 25316 4261 25344
rect 3384 25304 3390 25316
rect 4249 25313 4261 25316
rect 4295 25313 4307 25347
rect 5258 25344 5264 25356
rect 4249 25307 4307 25313
rect 4356 25316 5264 25344
rect 4356 25276 4384 25316
rect 5258 25304 5264 25316
rect 5316 25304 5322 25356
rect 7098 25344 7104 25356
rect 7059 25316 7104 25344
rect 7098 25304 7104 25316
rect 7156 25304 7162 25356
rect 7239 25347 7297 25353
rect 7239 25313 7251 25347
rect 7285 25313 7297 25347
rect 7374 25344 7380 25356
rect 7335 25316 7380 25344
rect 7239 25307 7297 25313
rect 5166 25276 5172 25288
rect 2740 25248 4384 25276
rect 5127 25248 5172 25276
rect 2740 25236 2746 25248
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 7254 25276 7282 25307
rect 7374 25304 7380 25316
rect 7432 25304 7438 25356
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25344 7527 25347
rect 7834 25344 7840 25356
rect 7515 25316 7840 25344
rect 7515 25313 7527 25316
rect 7469 25307 7527 25313
rect 7834 25304 7840 25316
rect 7892 25304 7898 25356
rect 8128 25353 8156 25384
rect 9508 25384 11152 25412
rect 9508 25353 9536 25384
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 12268 25412 12296 25440
rect 12437 25415 12495 25421
rect 12437 25412 12449 25415
rect 12268 25384 12449 25412
rect 12437 25381 12449 25384
rect 12483 25381 12495 25415
rect 12437 25375 12495 25381
rect 12526 25372 12532 25424
rect 12584 25412 12590 25424
rect 12584 25384 12629 25412
rect 12584 25372 12590 25384
rect 13170 25372 13176 25424
rect 13228 25412 13234 25424
rect 13541 25415 13599 25421
rect 13541 25412 13553 25415
rect 13228 25384 13553 25412
rect 13228 25372 13234 25384
rect 13541 25381 13553 25384
rect 13587 25381 13599 25415
rect 13648 25412 13676 25452
rect 13722 25440 13728 25492
rect 13780 25480 13786 25492
rect 13817 25483 13875 25489
rect 13817 25480 13829 25483
rect 13780 25452 13829 25480
rect 13780 25440 13786 25452
rect 13817 25449 13829 25452
rect 13863 25449 13875 25483
rect 13817 25443 13875 25449
rect 13906 25440 13912 25492
rect 13964 25480 13970 25492
rect 20898 25480 20904 25492
rect 13964 25452 20904 25480
rect 13964 25440 13970 25452
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 23382 25480 23388 25492
rect 23343 25452 23388 25480
rect 23382 25440 23388 25452
rect 23440 25440 23446 25492
rect 26602 25480 26608 25492
rect 26563 25452 26608 25480
rect 26602 25440 26608 25452
rect 26660 25440 26666 25492
rect 15004 25415 15062 25421
rect 13648 25384 14780 25412
rect 13541 25375 13599 25381
rect 8113 25347 8171 25353
rect 8113 25313 8125 25347
rect 8159 25313 8171 25347
rect 8113 25307 8171 25313
rect 9493 25347 9551 25353
rect 9493 25313 9505 25347
rect 9539 25313 9551 25347
rect 9493 25307 9551 25313
rect 9858 25304 9864 25356
rect 9916 25344 9922 25356
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 9916 25316 10149 25344
rect 9916 25304 9922 25316
rect 10137 25313 10149 25316
rect 10183 25313 10195 25347
rect 10137 25307 10195 25313
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25313 10931 25347
rect 10873 25307 10931 25313
rect 8018 25276 8024 25288
rect 7254 25248 8024 25276
rect 8018 25236 8024 25248
rect 8076 25236 8082 25288
rect 10888 25276 10916 25307
rect 10962 25304 10968 25356
rect 11020 25344 11026 25356
rect 11057 25347 11115 25353
rect 11057 25344 11069 25347
rect 11020 25316 11069 25344
rect 11020 25304 11026 25316
rect 11057 25313 11069 25316
rect 11103 25313 11115 25347
rect 11238 25344 11244 25356
rect 11199 25316 11244 25344
rect 11057 25307 11115 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 12250 25344 12256 25356
rect 12211 25316 12256 25344
rect 12250 25304 12256 25316
rect 12308 25304 12314 25356
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12802 25344 12808 25356
rect 12667 25316 12808 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 13265 25347 13323 25353
rect 13265 25313 13277 25347
rect 13311 25313 13323 25347
rect 13446 25344 13452 25356
rect 13407 25316 13452 25344
rect 13265 25307 13323 25313
rect 12066 25276 12072 25288
rect 10888 25248 12072 25276
rect 12066 25236 12072 25248
rect 12124 25236 12130 25288
rect 12710 25276 12716 25288
rect 12623 25248 12716 25276
rect 8573 25211 8631 25217
rect 8573 25177 8585 25211
rect 8619 25208 8631 25211
rect 10042 25208 10048 25220
rect 8619 25180 10048 25208
rect 8619 25177 8631 25180
rect 8573 25171 8631 25177
rect 10042 25168 10048 25180
rect 10100 25168 10106 25220
rect 11882 25168 11888 25220
rect 11940 25208 11946 25220
rect 12636 25208 12664 25248
rect 12710 25236 12716 25248
rect 12768 25276 12774 25288
rect 13078 25276 13084 25288
rect 12768 25248 13084 25276
rect 12768 25236 12774 25248
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13280 25276 13308 25307
rect 13446 25304 13452 25316
rect 13504 25304 13510 25356
rect 13633 25347 13691 25353
rect 13633 25313 13645 25347
rect 13679 25344 13691 25347
rect 13722 25344 13728 25356
rect 13679 25316 13728 25344
rect 13679 25313 13691 25316
rect 13633 25307 13691 25313
rect 13722 25304 13728 25316
rect 13780 25304 13786 25356
rect 14752 25353 14780 25384
rect 15004 25381 15016 25415
rect 15050 25412 15062 25415
rect 15194 25412 15200 25424
rect 15050 25384 15200 25412
rect 15050 25381 15062 25384
rect 15004 25375 15062 25381
rect 15194 25372 15200 25384
rect 15252 25372 15258 25424
rect 23109 25415 23167 25421
rect 23109 25381 23121 25415
rect 23155 25412 23167 25415
rect 23290 25412 23296 25424
rect 23155 25384 23296 25412
rect 23155 25381 23167 25384
rect 23109 25375 23167 25381
rect 23290 25372 23296 25384
rect 23348 25412 23354 25424
rect 24946 25412 24952 25424
rect 23348 25384 24952 25412
rect 23348 25372 23354 25384
rect 24946 25372 24952 25384
rect 25004 25372 25010 25424
rect 25222 25372 25228 25424
rect 25280 25412 25286 25424
rect 25470 25415 25528 25421
rect 25470 25412 25482 25415
rect 25280 25384 25482 25412
rect 25280 25372 25286 25384
rect 25470 25381 25482 25384
rect 25516 25381 25528 25415
rect 25470 25375 25528 25381
rect 14737 25347 14795 25353
rect 14737 25313 14749 25347
rect 14783 25313 14795 25347
rect 16666 25344 16672 25356
rect 16627 25316 16672 25344
rect 14737 25307 14795 25313
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 17310 25344 17316 25356
rect 17271 25316 17316 25344
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 17773 25347 17831 25353
rect 17773 25313 17785 25347
rect 17819 25313 17831 25347
rect 18138 25344 18144 25356
rect 18099 25316 18144 25344
rect 17773 25307 17831 25313
rect 13354 25276 13360 25288
rect 13267 25248 13360 25276
rect 13280 25208 13308 25248
rect 13354 25236 13360 25248
rect 13412 25276 13418 25288
rect 16761 25279 16819 25285
rect 13412 25248 13915 25276
rect 13412 25236 13418 25248
rect 11940 25180 12664 25208
rect 12728 25180 13308 25208
rect 11940 25168 11946 25180
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 2130 25140 2136 25152
rect 1627 25112 2136 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 2130 25100 2136 25112
rect 2188 25100 2194 25152
rect 4338 25140 4344 25152
rect 4299 25112 4344 25140
rect 4338 25100 4344 25112
rect 4396 25100 4402 25152
rect 7650 25140 7656 25152
rect 7611 25112 7656 25140
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 8202 25140 8208 25152
rect 8163 25112 8208 25140
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 9585 25143 9643 25149
rect 9585 25109 9597 25143
rect 9631 25140 9643 25143
rect 10134 25140 10140 25152
rect 9631 25112 10140 25140
rect 9631 25109 9643 25112
rect 9585 25103 9643 25109
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 10229 25143 10287 25149
rect 10229 25109 10241 25143
rect 10275 25140 10287 25143
rect 10594 25140 10600 25152
rect 10275 25112 10600 25140
rect 10275 25109 10287 25112
rect 10229 25103 10287 25109
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 12250 25100 12256 25152
rect 12308 25140 12314 25152
rect 12728 25140 12756 25180
rect 12308 25112 12756 25140
rect 12308 25100 12314 25112
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 13722 25140 13728 25152
rect 12860 25112 13728 25140
rect 12860 25100 12866 25112
rect 13722 25100 13728 25112
rect 13780 25100 13786 25152
rect 13887 25140 13915 25248
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 17497 25279 17555 25285
rect 17497 25276 17509 25279
rect 16807 25248 17509 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 17497 25245 17509 25248
rect 17543 25245 17555 25279
rect 17497 25239 17555 25245
rect 17034 25168 17040 25220
rect 17092 25208 17098 25220
rect 17788 25208 17816 25307
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 18325 25347 18383 25353
rect 18325 25313 18337 25347
rect 18371 25313 18383 25347
rect 18782 25344 18788 25356
rect 18743 25316 18788 25344
rect 18325 25307 18383 25313
rect 18340 25276 18368 25307
rect 18782 25304 18788 25316
rect 18840 25304 18846 25356
rect 22186 25304 22192 25356
rect 22244 25344 22250 25356
rect 22833 25347 22891 25353
rect 22833 25344 22845 25347
rect 22244 25316 22845 25344
rect 22244 25304 22250 25316
rect 22833 25313 22845 25316
rect 22879 25313 22891 25347
rect 22833 25307 22891 25313
rect 23017 25347 23075 25353
rect 23017 25313 23029 25347
rect 23063 25313 23075 25347
rect 23017 25307 23075 25313
rect 23201 25347 23259 25353
rect 23201 25313 23213 25347
rect 23247 25344 23259 25347
rect 24210 25344 24216 25356
rect 23247 25316 24216 25344
rect 23247 25313 23259 25316
rect 23201 25307 23259 25313
rect 18690 25276 18696 25288
rect 18340 25248 18696 25276
rect 18690 25236 18696 25248
rect 18748 25236 18754 25288
rect 23032 25276 23060 25307
rect 24210 25304 24216 25316
rect 24268 25304 24274 25356
rect 26050 25344 26056 25356
rect 25240 25316 26056 25344
rect 24762 25276 24768 25288
rect 23032 25248 24768 25276
rect 24762 25236 24768 25248
rect 24820 25236 24826 25288
rect 25240 25285 25268 25316
rect 26050 25304 26056 25316
rect 26108 25304 26114 25356
rect 27065 25347 27123 25353
rect 27065 25313 27077 25347
rect 27111 25344 27123 25347
rect 27154 25344 27160 25356
rect 27111 25316 27160 25344
rect 27111 25313 27123 25316
rect 27065 25307 27123 25313
rect 27154 25304 27160 25316
rect 27212 25304 27218 25356
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25245 25283 25279
rect 25225 25239 25283 25245
rect 17092 25180 17816 25208
rect 17865 25211 17923 25217
rect 17092 25168 17098 25180
rect 17865 25177 17877 25211
rect 17911 25208 17923 25211
rect 21818 25208 21824 25220
rect 17911 25180 21824 25208
rect 17911 25177 17923 25180
rect 17865 25171 17923 25177
rect 21818 25168 21824 25180
rect 21876 25168 21882 25220
rect 15102 25140 15108 25152
rect 13887 25112 15108 25140
rect 15102 25100 15108 25112
rect 15160 25100 15166 25152
rect 16114 25140 16120 25152
rect 16075 25112 16120 25140
rect 16114 25100 16120 25112
rect 16172 25100 16178 25152
rect 18322 25100 18328 25152
rect 18380 25140 18386 25152
rect 18877 25143 18935 25149
rect 18877 25140 18889 25143
rect 18380 25112 18889 25140
rect 18380 25100 18386 25112
rect 18877 25109 18889 25112
rect 18923 25109 18935 25143
rect 18877 25103 18935 25109
rect 1104 25050 28428 25072
rect 1104 24998 5536 25050
rect 5588 24998 5600 25050
rect 5652 24998 5664 25050
rect 5716 24998 5728 25050
rect 5780 24998 14644 25050
rect 14696 24998 14708 25050
rect 14760 24998 14772 25050
rect 14824 24998 14836 25050
rect 14888 24998 23752 25050
rect 23804 24998 23816 25050
rect 23868 24998 23880 25050
rect 23932 24998 23944 25050
rect 23996 24998 28428 25050
rect 1104 24976 28428 24998
rect 4338 24896 4344 24948
rect 4396 24936 4402 24948
rect 4396 24908 14412 24936
rect 4396 24896 4402 24908
rect 5258 24828 5264 24880
rect 5316 24868 5322 24880
rect 5353 24871 5411 24877
rect 5353 24868 5365 24871
rect 5316 24840 5365 24868
rect 5316 24828 5322 24840
rect 5353 24837 5365 24840
rect 5399 24837 5411 24871
rect 5353 24831 5411 24837
rect 7098 24828 7104 24880
rect 7156 24868 7162 24880
rect 7193 24871 7251 24877
rect 7193 24868 7205 24871
rect 7156 24840 7205 24868
rect 7156 24828 7162 24840
rect 7193 24837 7205 24840
rect 7239 24837 7251 24871
rect 7193 24831 7251 24837
rect 11422 24828 11428 24880
rect 11480 24868 11486 24880
rect 12066 24868 12072 24880
rect 11480 24840 12072 24868
rect 11480 24828 11486 24840
rect 12066 24828 12072 24840
rect 12124 24868 12130 24880
rect 12618 24868 12624 24880
rect 12124 24840 12624 24868
rect 12124 24828 12130 24840
rect 12618 24828 12624 24840
rect 12676 24828 12682 24880
rect 13265 24871 13323 24877
rect 13265 24837 13277 24871
rect 13311 24868 13323 24871
rect 13906 24868 13912 24880
rect 13311 24840 13912 24868
rect 13311 24837 13323 24840
rect 13265 24831 13323 24837
rect 13906 24828 13912 24840
rect 13964 24828 13970 24880
rect 2498 24800 2504 24812
rect 2240 24772 2504 24800
rect 1486 24692 1492 24744
rect 1544 24732 1550 24744
rect 2240 24741 2268 24772
rect 2498 24760 2504 24772
rect 2556 24800 2562 24812
rect 2682 24800 2688 24812
rect 2556 24772 2688 24800
rect 2556 24760 2562 24772
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 2866 24760 2872 24812
rect 2924 24800 2930 24812
rect 2924 24772 3280 24800
rect 2924 24760 2930 24772
rect 2225 24735 2283 24741
rect 1544 24704 1716 24732
rect 1544 24692 1550 24704
rect 1578 24664 1584 24676
rect 1539 24636 1584 24664
rect 1578 24624 1584 24636
rect 1636 24624 1642 24676
rect 1688 24664 1716 24704
rect 2225 24701 2237 24735
rect 2271 24701 2283 24735
rect 2225 24695 2283 24701
rect 2593 24735 2651 24741
rect 2593 24701 2605 24735
rect 2639 24732 2651 24735
rect 3142 24732 3148 24744
rect 2639 24704 3148 24732
rect 2639 24701 2651 24704
rect 2593 24695 2651 24701
rect 3142 24692 3148 24704
rect 3200 24692 3206 24744
rect 3252 24741 3280 24772
rect 5166 24760 5172 24812
rect 5224 24800 5230 24812
rect 7653 24803 7711 24809
rect 7653 24800 7665 24803
rect 5224 24772 7665 24800
rect 5224 24760 5230 24772
rect 7653 24769 7665 24772
rect 7699 24769 7711 24803
rect 7653 24763 7711 24769
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 10686 24800 10692 24812
rect 10367 24772 10692 24800
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24800 10839 24803
rect 12713 24803 12771 24809
rect 12713 24800 12725 24803
rect 10827 24772 12725 24800
rect 10827 24769 10839 24772
rect 10781 24763 10839 24769
rect 12713 24769 12725 24772
rect 12759 24769 12771 24803
rect 13630 24800 13636 24812
rect 12713 24763 12771 24769
rect 12912 24772 13636 24800
rect 3237 24735 3295 24741
rect 3237 24701 3249 24735
rect 3283 24732 3295 24735
rect 5184 24732 5212 24760
rect 10042 24732 10048 24744
rect 3283 24704 5212 24732
rect 7852 24704 9168 24732
rect 10003 24704 10048 24732
rect 3283 24701 3295 24704
rect 3237 24695 3295 24701
rect 2409 24667 2467 24673
rect 2409 24664 2421 24667
rect 1688 24636 2421 24664
rect 2409 24633 2421 24636
rect 2455 24633 2467 24667
rect 2409 24627 2467 24633
rect 2501 24667 2559 24673
rect 2501 24633 2513 24667
rect 2547 24664 2559 24667
rect 3326 24664 3332 24676
rect 2547 24636 3332 24664
rect 2547 24633 2559 24636
rect 2501 24627 2559 24633
rect 3326 24624 3332 24636
rect 3384 24624 3390 24676
rect 3504 24667 3562 24673
rect 3504 24633 3516 24667
rect 3550 24664 3562 24667
rect 4798 24664 4804 24676
rect 3550 24636 4804 24664
rect 3550 24633 3562 24636
rect 3504 24627 3562 24633
rect 4798 24624 4804 24636
rect 4856 24624 4862 24676
rect 5169 24667 5227 24673
rect 5169 24633 5181 24667
rect 5215 24664 5227 24667
rect 7009 24667 7067 24673
rect 7009 24664 7021 24667
rect 5215 24636 7021 24664
rect 5215 24633 5227 24636
rect 5169 24627 5227 24633
rect 7009 24633 7021 24636
rect 7055 24664 7067 24667
rect 7852 24664 7880 24704
rect 7055 24636 7880 24664
rect 7055 24633 7067 24636
rect 7009 24627 7067 24633
rect 1670 24596 1676 24608
rect 1631 24568 1676 24596
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 2774 24556 2780 24608
rect 2832 24596 2838 24608
rect 2832 24568 2877 24596
rect 2832 24556 2838 24568
rect 4522 24556 4528 24608
rect 4580 24596 4586 24608
rect 4617 24599 4675 24605
rect 4617 24596 4629 24599
rect 4580 24568 4629 24596
rect 4580 24556 4586 24568
rect 4617 24565 4629 24568
rect 4663 24565 4675 24599
rect 7852 24596 7880 24636
rect 7920 24667 7978 24673
rect 7920 24633 7932 24667
rect 7966 24664 7978 24667
rect 8570 24664 8576 24676
rect 7966 24636 8576 24664
rect 7966 24633 7978 24636
rect 7920 24627 7978 24633
rect 8570 24624 8576 24636
rect 8628 24624 8634 24676
rect 8110 24596 8116 24608
rect 7852 24568 8116 24596
rect 4617 24559 4675 24565
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 9033 24599 9091 24605
rect 9033 24596 9045 24599
rect 8996 24568 9045 24596
rect 8996 24556 9002 24568
rect 9033 24565 9045 24568
rect 9079 24565 9091 24599
rect 9140 24596 9168 24704
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 10134 24692 10140 24744
rect 10192 24732 10198 24744
rect 10229 24735 10287 24741
rect 10229 24732 10241 24735
rect 10192 24704 10241 24732
rect 10192 24692 10198 24704
rect 10229 24701 10241 24704
rect 10275 24701 10287 24735
rect 10229 24695 10287 24701
rect 10413 24735 10471 24741
rect 10413 24701 10425 24735
rect 10459 24701 10471 24735
rect 10594 24732 10600 24744
rect 10555 24704 10600 24732
rect 10413 24695 10471 24701
rect 10428 24664 10456 24695
rect 10594 24692 10600 24704
rect 10652 24692 10658 24744
rect 11054 24692 11060 24744
rect 11112 24732 11118 24744
rect 12069 24735 12127 24741
rect 12069 24732 12081 24735
rect 11112 24704 12081 24732
rect 11112 24692 11118 24704
rect 12069 24701 12081 24704
rect 12115 24701 12127 24735
rect 12069 24695 12127 24701
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24732 12219 24735
rect 12912 24732 12940 24772
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13998 24800 14004 24812
rect 13959 24772 14004 24800
rect 13998 24760 14004 24772
rect 14056 24760 14062 24812
rect 14384 24800 14412 24908
rect 14844 24908 15608 24936
rect 14461 24871 14519 24877
rect 14461 24837 14473 24871
rect 14507 24868 14519 24871
rect 14844 24868 14872 24908
rect 14507 24840 14872 24868
rect 14507 24837 14519 24840
rect 14461 24831 14519 24837
rect 14918 24828 14924 24880
rect 14976 24868 14982 24880
rect 14976 24840 15424 24868
rect 14976 24828 14982 24840
rect 14384 24772 14596 24800
rect 12207 24704 12940 24732
rect 12989 24735 13047 24741
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12989 24701 13001 24735
rect 13035 24732 13047 24735
rect 13078 24732 13084 24744
rect 13035 24704 13084 24732
rect 13035 24701 13047 24704
rect 12989 24695 13047 24701
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13262 24732 13268 24744
rect 13223 24704 13268 24732
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 14182 24732 14188 24744
rect 14143 24704 14188 24732
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 14568 24741 14596 24772
rect 14553 24735 14611 24741
rect 14332 24704 14377 24732
rect 14332 24692 14338 24704
rect 14553 24701 14565 24735
rect 14599 24701 14611 24735
rect 15286 24732 15292 24744
rect 15247 24704 15292 24732
rect 14553 24695 14611 24701
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 15396 24741 15424 24840
rect 15580 24812 15608 24908
rect 15654 24896 15660 24948
rect 15712 24936 15718 24948
rect 15712 24908 18180 24936
rect 15712 24896 15718 24908
rect 18049 24871 18107 24877
rect 18049 24837 18061 24871
rect 18095 24837 18107 24871
rect 18152 24868 18180 24908
rect 18690 24896 18696 24948
rect 18748 24936 18754 24948
rect 18877 24939 18935 24945
rect 18877 24936 18889 24939
rect 18748 24908 18889 24936
rect 18748 24896 18754 24908
rect 18877 24905 18889 24908
rect 18923 24905 18935 24939
rect 18877 24899 18935 24905
rect 19058 24868 19064 24880
rect 18152 24840 19064 24868
rect 18049 24831 18107 24837
rect 15562 24800 15568 24812
rect 15523 24772 15568 24800
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 16301 24803 16359 24809
rect 16301 24769 16313 24803
rect 16347 24800 16359 24803
rect 17497 24803 17555 24809
rect 17497 24800 17509 24803
rect 16347 24772 17509 24800
rect 16347 24769 16359 24772
rect 16301 24763 16359 24769
rect 17497 24769 17509 24772
rect 17543 24769 17555 24803
rect 18064 24800 18092 24831
rect 19058 24828 19064 24840
rect 19116 24868 19122 24880
rect 22094 24868 22100 24880
rect 19116 24840 22100 24868
rect 19116 24828 19122 24840
rect 22094 24828 22100 24840
rect 22152 24828 22158 24880
rect 23569 24871 23627 24877
rect 23569 24837 23581 24871
rect 23615 24837 23627 24871
rect 23569 24831 23627 24837
rect 18064 24772 22094 24800
rect 17497 24763 17555 24769
rect 15381 24735 15439 24741
rect 15381 24701 15393 24735
rect 15427 24701 15439 24735
rect 15654 24732 15660 24744
rect 15615 24704 15660 24732
rect 15381 24695 15439 24701
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 16206 24732 16212 24744
rect 16167 24704 16212 24732
rect 16206 24692 16212 24704
rect 16264 24692 16270 24744
rect 17313 24735 17371 24741
rect 17313 24701 17325 24735
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 10778 24664 10784 24676
rect 10428 24636 10784 24664
rect 10778 24624 10784 24636
rect 10836 24624 10842 24676
rect 13538 24664 13544 24676
rect 13499 24636 13544 24664
rect 13538 24624 13544 24636
rect 13596 24624 13602 24676
rect 15105 24667 15163 24673
rect 15105 24633 15117 24667
rect 15151 24664 15163 24667
rect 17328 24664 17356 24695
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 17773 24735 17831 24741
rect 17773 24732 17785 24735
rect 17460 24704 17785 24732
rect 17460 24692 17466 24704
rect 17773 24701 17785 24704
rect 17819 24701 17831 24735
rect 18138 24732 18144 24744
rect 18051 24704 18144 24732
rect 17773 24695 17831 24701
rect 18138 24692 18144 24704
rect 18196 24692 18202 24744
rect 18322 24732 18328 24744
rect 18283 24704 18328 24732
rect 18322 24692 18328 24704
rect 18380 24692 18386 24744
rect 18785 24735 18843 24741
rect 18785 24701 18797 24735
rect 18831 24732 18843 24735
rect 18874 24732 18880 24744
rect 18831 24704 18880 24732
rect 18831 24701 18843 24704
rect 18785 24695 18843 24701
rect 18874 24692 18880 24704
rect 18932 24692 18938 24744
rect 21177 24735 21235 24741
rect 21177 24701 21189 24735
rect 21223 24732 21235 24735
rect 21450 24732 21456 24744
rect 21223 24704 21456 24732
rect 21223 24701 21235 24704
rect 21177 24695 21235 24701
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 22066 24732 22094 24772
rect 23017 24735 23075 24741
rect 23017 24732 23029 24735
rect 22066 24704 23029 24732
rect 23017 24701 23029 24704
rect 23063 24701 23075 24735
rect 23198 24732 23204 24744
rect 23159 24704 23204 24732
rect 23017 24695 23075 24701
rect 23198 24692 23204 24704
rect 23256 24692 23262 24744
rect 23382 24732 23388 24744
rect 23343 24704 23388 24732
rect 23382 24692 23388 24704
rect 23440 24692 23446 24744
rect 15151 24636 17356 24664
rect 18156 24664 18184 24692
rect 18966 24664 18972 24676
rect 18156 24636 18972 24664
rect 15151 24633 15163 24636
rect 15105 24627 15163 24633
rect 18966 24624 18972 24636
rect 19024 24624 19030 24676
rect 21082 24624 21088 24676
rect 21140 24664 21146 24676
rect 23216 24664 23244 24692
rect 21140 24636 23244 24664
rect 21140 24624 21146 24636
rect 23290 24624 23296 24676
rect 23348 24664 23354 24676
rect 23584 24664 23612 24831
rect 24029 24735 24087 24741
rect 24029 24701 24041 24735
rect 24075 24732 24087 24735
rect 24118 24732 24124 24744
rect 24075 24704 24124 24732
rect 24075 24701 24087 24704
rect 24029 24695 24087 24701
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 26142 24732 26148 24744
rect 26103 24704 26148 24732
rect 26142 24692 26148 24704
rect 26200 24692 26206 24744
rect 26513 24735 26571 24741
rect 26513 24701 26525 24735
rect 26559 24732 26571 24735
rect 26602 24732 26608 24744
rect 26559 24704 26608 24732
rect 26559 24701 26571 24704
rect 26513 24695 26571 24701
rect 26602 24692 26608 24704
rect 26660 24692 26666 24744
rect 24274 24667 24332 24673
rect 24274 24664 24286 24667
rect 23348 24636 23393 24664
rect 23584 24636 24286 24664
rect 23348 24624 23354 24636
rect 24274 24633 24286 24636
rect 24320 24633 24332 24667
rect 26326 24664 26332 24676
rect 26287 24636 26332 24664
rect 24274 24627 24332 24633
rect 26326 24624 26332 24636
rect 26384 24624 26390 24676
rect 26418 24624 26424 24676
rect 26476 24664 26482 24676
rect 26476 24636 26521 24664
rect 26476 24624 26482 24636
rect 17494 24596 17500 24608
rect 9140 24568 17500 24596
rect 9033 24559 9091 24565
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 21269 24599 21327 24605
rect 21269 24565 21281 24599
rect 21315 24596 21327 24599
rect 22922 24596 22928 24608
rect 21315 24568 22928 24596
rect 21315 24565 21327 24568
rect 21269 24559 21327 24565
rect 22922 24556 22928 24568
rect 22980 24556 22986 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 25409 24599 25467 24605
rect 25409 24596 25421 24599
rect 23440 24568 25421 24596
rect 23440 24556 23446 24568
rect 25409 24565 25421 24568
rect 25455 24596 25467 24599
rect 26234 24596 26240 24608
rect 25455 24568 26240 24596
rect 25455 24565 25467 24568
rect 25409 24559 25467 24565
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 26694 24596 26700 24608
rect 26655 24568 26700 24596
rect 26694 24556 26700 24568
rect 26752 24556 26758 24608
rect 1104 24506 28428 24528
rect 1104 24454 10090 24506
rect 10142 24454 10154 24506
rect 10206 24454 10218 24506
rect 10270 24454 10282 24506
rect 10334 24454 19198 24506
rect 19250 24454 19262 24506
rect 19314 24454 19326 24506
rect 19378 24454 19390 24506
rect 19442 24454 28428 24506
rect 1104 24432 28428 24454
rect 3326 24392 3332 24404
rect 3287 24364 3332 24392
rect 3326 24352 3332 24364
rect 3384 24352 3390 24404
rect 4798 24392 4804 24404
rect 3436 24364 4660 24392
rect 4759 24364 4804 24392
rect 2216 24327 2274 24333
rect 2216 24293 2228 24327
rect 2262 24324 2274 24327
rect 2774 24324 2780 24336
rect 2262 24296 2780 24324
rect 2262 24293 2274 24296
rect 2216 24287 2274 24293
rect 2774 24284 2780 24296
rect 2832 24284 2838 24336
rect 2866 24284 2872 24336
rect 2924 24284 2930 24336
rect 3142 24284 3148 24336
rect 3200 24324 3206 24336
rect 3436 24324 3464 24364
rect 4522 24324 4528 24336
rect 3200 24296 3464 24324
rect 4483 24296 4528 24324
rect 3200 24284 3206 24296
rect 4522 24284 4528 24296
rect 4580 24284 4586 24336
rect 4632 24324 4660 24364
rect 4798 24352 4804 24364
rect 4856 24352 4862 24404
rect 7558 24392 7564 24404
rect 6012 24364 7564 24392
rect 5537 24327 5595 24333
rect 5537 24324 5549 24327
rect 4632 24296 5549 24324
rect 1949 24259 2007 24265
rect 1949 24225 1961 24259
rect 1995 24256 2007 24259
rect 2884 24256 2912 24284
rect 1995 24228 2912 24256
rect 4249 24259 4307 24265
rect 1995 24225 2007 24228
rect 1949 24219 2007 24225
rect 4249 24225 4261 24259
rect 4295 24225 4307 24259
rect 4430 24256 4436 24268
rect 4391 24228 4436 24256
rect 4249 24219 4307 24225
rect 4264 24188 4292 24219
rect 4430 24216 4436 24228
rect 4488 24216 4494 24268
rect 4632 24265 4660 24296
rect 5537 24293 5549 24296
rect 5583 24324 5595 24327
rect 5902 24324 5908 24336
rect 5583 24296 5908 24324
rect 5583 24293 5595 24296
rect 5537 24287 5595 24293
rect 5902 24284 5908 24296
rect 5960 24284 5966 24336
rect 4617 24259 4675 24265
rect 4617 24225 4629 24259
rect 4663 24225 4675 24259
rect 4617 24219 4675 24225
rect 5353 24259 5411 24265
rect 5353 24225 5365 24259
rect 5399 24256 5411 24259
rect 6012 24256 6040 24364
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 8570 24392 8576 24404
rect 8531 24364 8576 24392
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 13173 24395 13231 24401
rect 13173 24361 13185 24395
rect 13219 24392 13231 24395
rect 13538 24392 13544 24404
rect 13219 24364 13544 24392
rect 13219 24361 13231 24364
rect 13173 24355 13231 24361
rect 13538 24352 13544 24364
rect 13596 24352 13602 24404
rect 15194 24352 15200 24404
rect 15252 24392 15258 24404
rect 15289 24395 15347 24401
rect 15289 24392 15301 24395
rect 15252 24364 15301 24392
rect 15252 24352 15258 24364
rect 15289 24361 15301 24364
rect 15335 24361 15347 24395
rect 15289 24355 15347 24361
rect 15930 24352 15936 24404
rect 15988 24392 15994 24404
rect 22646 24392 22652 24404
rect 15988 24364 22652 24392
rect 15988 24352 15994 24364
rect 22646 24352 22652 24364
rect 22704 24392 22710 24404
rect 26418 24392 26424 24404
rect 22704 24364 23060 24392
rect 22704 24352 22710 24364
rect 6356 24327 6414 24333
rect 6356 24293 6368 24327
rect 6402 24324 6414 24327
rect 7650 24324 7656 24336
rect 6402 24296 7656 24324
rect 6402 24293 6414 24296
rect 6356 24287 6414 24293
rect 7650 24284 7656 24296
rect 7708 24284 7714 24336
rect 8297 24327 8355 24333
rect 8297 24293 8309 24327
rect 8343 24324 8355 24327
rect 8938 24324 8944 24336
rect 8343 24296 8944 24324
rect 8343 24293 8355 24296
rect 8297 24287 8355 24293
rect 8938 24284 8944 24296
rect 8996 24284 9002 24336
rect 14366 24284 14372 24336
rect 14424 24324 14430 24336
rect 14921 24327 14979 24333
rect 14921 24324 14933 24327
rect 14424 24296 14933 24324
rect 14424 24284 14430 24296
rect 14921 24293 14933 24296
rect 14967 24293 14979 24327
rect 14921 24287 14979 24293
rect 15013 24327 15071 24333
rect 15013 24293 15025 24327
rect 15059 24324 15071 24327
rect 17494 24324 17500 24336
rect 15059 24296 15792 24324
rect 17455 24296 17500 24324
rect 15059 24293 15071 24296
rect 15013 24287 15071 24293
rect 5399 24228 6040 24256
rect 5399 24225 5411 24228
rect 5353 24219 5411 24225
rect 7098 24216 7104 24268
rect 7156 24256 7162 24268
rect 8021 24259 8079 24265
rect 8021 24256 8033 24259
rect 7156 24228 8033 24256
rect 7156 24216 7162 24228
rect 8021 24225 8033 24228
rect 8067 24225 8079 24259
rect 8021 24219 8079 24225
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24225 8263 24259
rect 8389 24259 8447 24265
rect 8389 24256 8401 24259
rect 8205 24219 8263 24225
rect 8312 24228 8401 24256
rect 5258 24188 5264 24200
rect 4264 24160 5264 24188
rect 5258 24148 5264 24160
rect 5316 24148 5322 24200
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24157 6147 24191
rect 6089 24151 6147 24157
rect 5166 24080 5172 24132
rect 5224 24120 5230 24132
rect 6104 24120 6132 24151
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 8220 24188 8248 24219
rect 7708 24160 8248 24188
rect 7708 24148 7714 24160
rect 5224 24092 6132 24120
rect 5224 24080 5230 24092
rect 7834 24080 7840 24132
rect 7892 24120 7898 24132
rect 8312 24120 8340 24228
rect 8389 24225 8401 24228
rect 8435 24225 8447 24259
rect 8389 24219 8447 24225
rect 9490 24216 9496 24268
rect 9548 24256 9554 24268
rect 9861 24259 9919 24265
rect 9861 24256 9873 24259
rect 9548 24228 9873 24256
rect 9548 24216 9554 24228
rect 9861 24225 9873 24228
rect 9907 24225 9919 24259
rect 9861 24219 9919 24225
rect 9950 24216 9956 24268
rect 10008 24256 10014 24268
rect 10117 24259 10175 24265
rect 10117 24256 10129 24259
rect 10008 24228 10129 24256
rect 10008 24216 10014 24228
rect 10117 24225 10129 24228
rect 10163 24225 10175 24259
rect 10117 24219 10175 24225
rect 13081 24259 13139 24265
rect 13081 24225 13093 24259
rect 13127 24256 13139 24259
rect 13170 24256 13176 24268
rect 13127 24228 13176 24256
rect 13127 24225 13139 24228
rect 13081 24219 13139 24225
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 14737 24259 14795 24265
rect 14737 24225 14749 24259
rect 14783 24225 14795 24259
rect 14737 24219 14795 24225
rect 15105 24259 15163 24265
rect 15105 24225 15117 24259
rect 15151 24256 15163 24259
rect 15470 24256 15476 24268
rect 15151 24228 15476 24256
rect 15151 24225 15163 24228
rect 15105 24219 15163 24225
rect 14752 24188 14780 24219
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 15764 24265 15792 24296
rect 17494 24284 17500 24296
rect 17552 24284 17558 24336
rect 22741 24327 22799 24333
rect 22741 24324 22753 24327
rect 21284 24296 22753 24324
rect 15749 24259 15807 24265
rect 15749 24225 15761 24259
rect 15795 24256 15807 24259
rect 16114 24256 16120 24268
rect 15795 24228 16120 24256
rect 15795 24225 15807 24228
rect 15749 24219 15807 24225
rect 16114 24216 16120 24228
rect 16172 24216 16178 24268
rect 19518 24216 19524 24268
rect 19576 24256 19582 24268
rect 21284 24265 21312 24296
rect 22741 24293 22753 24296
rect 22787 24293 22799 24327
rect 22741 24287 22799 24293
rect 20533 24259 20591 24265
rect 20533 24256 20545 24259
rect 19576 24228 20545 24256
rect 19576 24216 19582 24228
rect 20533 24225 20545 24228
rect 20579 24225 20591 24259
rect 20533 24219 20591 24225
rect 21269 24259 21327 24265
rect 21269 24225 21281 24259
rect 21315 24225 21327 24259
rect 21269 24219 21327 24225
rect 21729 24259 21787 24265
rect 21729 24225 21741 24259
rect 21775 24225 21787 24259
rect 21729 24219 21787 24225
rect 15194 24188 15200 24200
rect 14752 24160 15200 24188
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 15286 24148 15292 24200
rect 15344 24188 15350 24200
rect 15841 24191 15899 24197
rect 15841 24188 15853 24191
rect 15344 24160 15853 24188
rect 15344 24148 15350 24160
rect 15841 24157 15853 24160
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 20625 24191 20683 24197
rect 20625 24157 20637 24191
rect 20671 24188 20683 24191
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 20671 24160 21465 24188
rect 20671 24157 20683 24160
rect 20625 24151 20683 24157
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 7892 24092 8340 24120
rect 7892 24080 7898 24092
rect 12802 24080 12808 24132
rect 12860 24120 12866 24132
rect 12986 24120 12992 24132
rect 12860 24092 12992 24120
rect 12860 24080 12866 24092
rect 12986 24080 12992 24092
rect 13044 24080 13050 24132
rect 13906 24080 13912 24132
rect 13964 24120 13970 24132
rect 17402 24120 17408 24132
rect 13964 24092 17408 24120
rect 13964 24080 13970 24092
rect 17402 24080 17408 24092
rect 17460 24080 17466 24132
rect 17678 24120 17684 24132
rect 17639 24092 17684 24120
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 7466 24052 7472 24064
rect 7427 24024 7472 24052
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 11241 24055 11299 24061
rect 11241 24052 11253 24055
rect 9732 24024 11253 24052
rect 9732 24012 9738 24024
rect 11241 24021 11253 24024
rect 11287 24021 11299 24055
rect 11241 24015 11299 24021
rect 13998 24012 14004 24064
rect 14056 24052 14062 24064
rect 16206 24052 16212 24064
rect 14056 24024 16212 24052
rect 14056 24012 14062 24024
rect 16206 24012 16212 24024
rect 16264 24012 16270 24064
rect 17420 24052 17448 24080
rect 21744 24052 21772 24219
rect 22094 24216 22100 24268
rect 22152 24256 22158 24268
rect 22281 24259 22339 24265
rect 22152 24228 22197 24256
rect 22152 24216 22158 24228
rect 22281 24225 22293 24259
rect 22327 24256 22339 24259
rect 22462 24256 22468 24268
rect 22327 24228 22468 24256
rect 22327 24225 22339 24228
rect 22281 24219 22339 24225
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 22922 24256 22928 24268
rect 22883 24228 22928 24256
rect 22922 24216 22928 24228
rect 22980 24216 22986 24268
rect 23032 24265 23060 24364
rect 25608 24364 26424 24392
rect 25501 24327 25559 24333
rect 25501 24324 25513 24327
rect 23308 24296 25513 24324
rect 23308 24265 23336 24296
rect 25501 24293 25513 24296
rect 25547 24293 25559 24327
rect 25501 24287 25559 24293
rect 23017 24259 23075 24265
rect 23017 24225 23029 24259
rect 23063 24225 23075 24259
rect 23017 24219 23075 24225
rect 23293 24259 23351 24265
rect 23293 24225 23305 24259
rect 23339 24225 23351 24259
rect 23293 24219 23351 24225
rect 25409 24259 25467 24265
rect 25409 24225 25421 24259
rect 25455 24256 25467 24259
rect 25608 24256 25636 24364
rect 26418 24352 26424 24364
rect 26476 24392 26482 24404
rect 27433 24395 27491 24401
rect 27433 24392 27445 24395
rect 26476 24364 27445 24392
rect 26476 24352 26482 24364
rect 27433 24361 27445 24364
rect 27479 24361 27491 24395
rect 27433 24355 27491 24361
rect 26320 24327 26378 24333
rect 26320 24293 26332 24327
rect 26366 24324 26378 24327
rect 26694 24324 26700 24336
rect 26366 24296 26700 24324
rect 26366 24293 26378 24296
rect 26320 24287 26378 24293
rect 26694 24284 26700 24296
rect 26752 24284 26758 24336
rect 25455 24228 25636 24256
rect 25455 24225 25467 24228
rect 25409 24219 25467 24225
rect 26050 24188 26056 24200
rect 26011 24160 26056 24188
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 22005 24123 22063 24129
rect 22005 24089 22017 24123
rect 22051 24120 22063 24123
rect 22094 24120 22100 24132
rect 22051 24092 22100 24120
rect 22051 24089 22063 24092
rect 22005 24083 22063 24089
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 22186 24052 22192 24064
rect 17420 24024 22192 24052
rect 22186 24012 22192 24024
rect 22244 24012 22250 24064
rect 23014 24012 23020 24064
rect 23072 24052 23078 24064
rect 23201 24055 23259 24061
rect 23201 24052 23213 24055
rect 23072 24024 23213 24052
rect 23072 24012 23078 24024
rect 23201 24021 23213 24024
rect 23247 24021 23259 24055
rect 23201 24015 23259 24021
rect 1104 23962 28428 23984
rect 1104 23910 5536 23962
rect 5588 23910 5600 23962
rect 5652 23910 5664 23962
rect 5716 23910 5728 23962
rect 5780 23910 14644 23962
rect 14696 23910 14708 23962
rect 14760 23910 14772 23962
rect 14824 23910 14836 23962
rect 14888 23910 23752 23962
rect 23804 23910 23816 23962
rect 23868 23910 23880 23962
rect 23932 23910 23944 23962
rect 23996 23910 28428 23962
rect 1104 23888 28428 23910
rect 2866 23848 2872 23860
rect 2516 23820 2872 23848
rect 2516 23721 2544 23820
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 5721 23851 5779 23857
rect 5721 23817 5733 23851
rect 5767 23848 5779 23851
rect 6914 23848 6920 23860
rect 5767 23820 6920 23848
rect 5767 23817 5779 23820
rect 5721 23811 5779 23817
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 7558 23808 7564 23860
rect 7616 23848 7622 23860
rect 7616 23820 17448 23848
rect 7616 23808 7622 23820
rect 4893 23783 4951 23789
rect 4893 23749 4905 23783
rect 4939 23780 4951 23783
rect 9950 23780 9956 23792
rect 4939 23752 9674 23780
rect 9911 23752 9956 23780
rect 4939 23749 4951 23752
rect 4893 23743 4951 23749
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23681 2559 23715
rect 7834 23712 7840 23724
rect 7795 23684 7840 23712
rect 2501 23675 2559 23681
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 9646 23712 9674 23752
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 16206 23780 16212 23792
rect 10051 23752 16212 23780
rect 10051 23712 10079 23752
rect 16206 23740 16212 23752
rect 16264 23740 16270 23792
rect 10502 23712 10508 23724
rect 9646 23684 10079 23712
rect 10268 23684 10508 23712
rect 1578 23604 1584 23656
rect 1636 23644 1642 23656
rect 1765 23647 1823 23653
rect 1765 23644 1777 23647
rect 1636 23616 1777 23644
rect 1636 23604 1642 23616
rect 1765 23613 1777 23616
rect 1811 23613 1823 23647
rect 1765 23607 1823 23613
rect 1780 23508 1808 23607
rect 4522 23604 4528 23656
rect 4580 23644 4586 23656
rect 4801 23647 4859 23653
rect 4801 23644 4813 23647
rect 4580 23616 4813 23644
rect 4580 23604 4586 23616
rect 4801 23613 4813 23616
rect 4847 23613 4859 23647
rect 4801 23607 4859 23613
rect 5445 23647 5503 23653
rect 5445 23613 5457 23647
rect 5491 23644 5503 23647
rect 7466 23644 7472 23656
rect 5491 23616 7472 23644
rect 5491 23613 5503 23616
rect 5445 23607 5503 23613
rect 7466 23604 7472 23616
rect 7524 23604 7530 23656
rect 7558 23604 7564 23656
rect 7616 23644 7622 23656
rect 9398 23644 9404 23656
rect 7616 23616 7661 23644
rect 9359 23616 9404 23644
rect 7616 23604 7622 23616
rect 9398 23604 9404 23616
rect 9456 23604 9462 23656
rect 9674 23644 9680 23656
rect 9508 23616 9680 23644
rect 2768 23579 2826 23585
rect 2768 23545 2780 23579
rect 2814 23576 2826 23579
rect 3050 23576 3056 23588
rect 2814 23548 3056 23576
rect 2814 23545 2826 23548
rect 2768 23539 2826 23545
rect 3050 23536 3056 23548
rect 3108 23536 3114 23588
rect 9508 23576 9536 23616
rect 9674 23604 9680 23616
rect 9732 23604 9738 23656
rect 9769 23647 9827 23653
rect 9769 23613 9781 23647
rect 9815 23644 9827 23647
rect 10268 23644 10296 23684
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10778 23712 10784 23724
rect 10691 23684 10784 23712
rect 10778 23672 10784 23684
rect 10836 23712 10842 23724
rect 11330 23712 11336 23724
rect 10836 23684 11336 23712
rect 10836 23672 10842 23684
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 13354 23672 13360 23724
rect 13412 23672 13418 23724
rect 13722 23712 13728 23724
rect 13464 23684 13728 23712
rect 10410 23644 10416 23656
rect 9815 23616 10296 23644
rect 10371 23616 10416 23644
rect 9815 23613 9827 23616
rect 9769 23607 9827 23613
rect 10410 23604 10416 23616
rect 10468 23604 10474 23656
rect 10594 23644 10600 23656
rect 10555 23616 10600 23644
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 10689 23647 10747 23653
rect 10689 23613 10701 23647
rect 10735 23644 10747 23647
rect 10962 23644 10968 23656
rect 10735 23616 10824 23644
rect 10923 23616 10968 23644
rect 10735 23613 10747 23616
rect 10689 23607 10747 23613
rect 10796 23588 10824 23616
rect 10962 23604 10968 23616
rect 11020 23604 11026 23656
rect 13081 23647 13139 23653
rect 13081 23613 13093 23647
rect 13127 23644 13139 23647
rect 13372 23644 13400 23672
rect 13464 23653 13492 23684
rect 13722 23672 13728 23684
rect 13780 23712 13786 23724
rect 15470 23712 15476 23724
rect 13780 23684 15476 23712
rect 13780 23672 13786 23684
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 13127 23616 13400 23644
rect 13449 23647 13507 23653
rect 13127 23613 13139 23616
rect 13081 23607 13139 23613
rect 13449 23613 13461 23647
rect 13495 23613 13507 23647
rect 14090 23644 14096 23656
rect 14051 23616 14096 23644
rect 13449 23607 13507 23613
rect 14090 23604 14096 23616
rect 14148 23604 14154 23656
rect 15194 23604 15200 23656
rect 15252 23644 15258 23656
rect 17420 23653 17448 23820
rect 17678 23808 17684 23860
rect 17736 23848 17742 23860
rect 19518 23848 19524 23860
rect 17736 23820 19104 23848
rect 19479 23820 19524 23848
rect 17736 23808 17742 23820
rect 19076 23780 19104 23820
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19628 23820 24992 23848
rect 19628 23780 19656 23820
rect 19076 23752 19656 23780
rect 23017 23783 23075 23789
rect 23017 23749 23029 23783
rect 23063 23780 23075 23783
rect 23198 23780 23204 23792
rect 23063 23752 23204 23780
rect 23063 23749 23075 23752
rect 23017 23743 23075 23749
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 22704 23684 22876 23712
rect 22704 23672 22710 23684
rect 16025 23647 16083 23653
rect 16025 23644 16037 23647
rect 15252 23616 16037 23644
rect 15252 23604 15258 23616
rect 16025 23613 16037 23616
rect 16071 23613 16083 23647
rect 16025 23607 16083 23613
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23644 18199 23647
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 18187 23616 20085 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 20073 23613 20085 23616
rect 20119 23613 20131 23647
rect 22738 23644 22744 23656
rect 22699 23616 22744 23644
rect 20073 23607 20131 23613
rect 3712 23548 9536 23576
rect 9585 23579 9643 23585
rect 3712 23508 3740 23548
rect 9585 23545 9597 23579
rect 9631 23545 9643 23579
rect 9585 23539 9643 23545
rect 3878 23508 3884 23520
rect 1780 23480 3740 23508
rect 3839 23480 3884 23508
rect 3878 23468 3884 23480
rect 3936 23468 3942 23520
rect 5905 23511 5963 23517
rect 5905 23477 5917 23511
rect 5951 23508 5963 23511
rect 6730 23508 6736 23520
rect 5951 23480 6736 23508
rect 5951 23477 5963 23480
rect 5905 23471 5963 23477
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 9600 23508 9628 23539
rect 10778 23536 10784 23588
rect 10836 23536 10842 23588
rect 13170 23576 13176 23588
rect 11072 23548 13176 23576
rect 11072 23508 11100 23548
rect 13170 23536 13176 23548
rect 13228 23576 13234 23588
rect 13265 23579 13323 23585
rect 13265 23576 13277 23579
rect 13228 23548 13277 23576
rect 13228 23536 13234 23548
rect 13265 23545 13277 23548
rect 13311 23545 13323 23579
rect 13265 23539 13323 23545
rect 13357 23579 13415 23585
rect 13357 23545 13369 23579
rect 13403 23576 13415 23579
rect 14108 23576 14136 23604
rect 15286 23576 15292 23588
rect 13403 23548 14136 23576
rect 15247 23548 15292 23576
rect 13403 23545 13415 23548
rect 13357 23539 13415 23545
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 17218 23536 17224 23588
rect 17276 23576 17282 23588
rect 18156 23576 18184 23607
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 22848 23653 22876 23684
rect 22848 23647 22921 23653
rect 22848 23616 22875 23647
rect 22863 23613 22875 23616
rect 22909 23613 22921 23647
rect 22863 23607 22921 23613
rect 23109 23647 23167 23653
rect 23109 23613 23121 23647
rect 23155 23613 23167 23647
rect 23934 23644 23940 23656
rect 23895 23616 23940 23644
rect 23109 23607 23167 23613
rect 18414 23585 18420 23588
rect 17276 23548 18184 23576
rect 17276 23536 17282 23548
rect 18408 23539 18420 23585
rect 18472 23576 18478 23588
rect 20340 23579 20398 23585
rect 18472 23548 18508 23576
rect 18414 23536 18420 23539
rect 18472 23536 18478 23548
rect 20340 23545 20352 23579
rect 20386 23576 20398 23579
rect 20622 23576 20628 23588
rect 20386 23548 20628 23576
rect 20386 23545 20398 23548
rect 20340 23539 20398 23545
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 21542 23536 21548 23588
rect 21600 23576 21606 23588
rect 23124 23576 23152 23607
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24964 23644 24992 23820
rect 26418 23672 26424 23724
rect 26476 23672 26482 23724
rect 26142 23644 26148 23656
rect 24964 23616 26148 23644
rect 26142 23604 26148 23616
rect 26200 23604 26206 23656
rect 26329 23647 26387 23653
rect 26329 23613 26341 23647
rect 26375 23644 26387 23647
rect 26436 23644 26464 23672
rect 26375 23616 26464 23644
rect 26513 23647 26571 23653
rect 26375 23613 26387 23616
rect 26329 23607 26387 23613
rect 26513 23613 26525 23647
rect 26559 23644 26571 23647
rect 26602 23644 26608 23656
rect 26559 23616 26608 23644
rect 26559 23613 26571 23616
rect 26513 23607 26571 23613
rect 26602 23604 26608 23616
rect 26660 23604 26666 23656
rect 24210 23585 24216 23588
rect 21600 23548 23152 23576
rect 21600 23536 21606 23548
rect 24204 23539 24216 23585
rect 24268 23576 24274 23588
rect 26421 23579 26479 23585
rect 24268 23548 24304 23576
rect 24210 23536 24216 23539
rect 24268 23536 24274 23548
rect 26421 23545 26433 23579
rect 26467 23545 26479 23579
rect 26421 23539 26479 23545
rect 9600 23480 11100 23508
rect 11149 23511 11207 23517
rect 11149 23477 11161 23511
rect 11195 23508 11207 23511
rect 12986 23508 12992 23520
rect 11195 23480 12992 23508
rect 11195 23477 11207 23480
rect 11149 23471 11207 23477
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 13630 23508 13636 23520
rect 13591 23480 13636 23508
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 14182 23508 14188 23520
rect 14143 23480 14188 23508
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 15010 23468 15016 23520
rect 15068 23508 15074 23520
rect 15381 23511 15439 23517
rect 15381 23508 15393 23511
rect 15068 23480 15393 23508
rect 15068 23468 15074 23480
rect 15381 23477 15393 23480
rect 15427 23477 15439 23511
rect 15381 23471 15439 23477
rect 15838 23468 15844 23520
rect 15896 23508 15902 23520
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 15896 23480 16129 23508
rect 15896 23468 15902 23480
rect 16117 23477 16129 23480
rect 16163 23477 16175 23511
rect 16117 23471 16175 23477
rect 17497 23511 17555 23517
rect 17497 23477 17509 23511
rect 17543 23508 17555 23511
rect 17954 23508 17960 23520
rect 17543 23480 17960 23508
rect 17543 23477 17555 23480
rect 17497 23471 17555 23477
rect 17954 23468 17960 23480
rect 18012 23508 18018 23520
rect 21266 23508 21272 23520
rect 18012 23480 21272 23508
rect 18012 23468 18018 23480
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 21450 23508 21456 23520
rect 21411 23480 21456 23508
rect 21450 23468 21456 23480
rect 21508 23468 21514 23520
rect 22557 23511 22615 23517
rect 22557 23477 22569 23511
rect 22603 23508 22615 23511
rect 23566 23508 23572 23520
rect 22603 23480 23572 23508
rect 22603 23477 22615 23480
rect 22557 23471 22615 23477
rect 23566 23468 23572 23480
rect 23624 23468 23630 23520
rect 25314 23468 25320 23520
rect 25372 23508 25378 23520
rect 25372 23480 25417 23508
rect 25372 23468 25378 23480
rect 26142 23468 26148 23520
rect 26200 23508 26206 23520
rect 26436 23508 26464 23539
rect 26694 23508 26700 23520
rect 26200 23480 26464 23508
rect 26655 23480 26700 23508
rect 26200 23468 26206 23480
rect 26694 23468 26700 23480
rect 26752 23468 26758 23520
rect 1104 23418 28428 23440
rect 1104 23366 10090 23418
rect 10142 23366 10154 23418
rect 10206 23366 10218 23418
rect 10270 23366 10282 23418
rect 10334 23366 19198 23418
rect 19250 23366 19262 23418
rect 19314 23366 19326 23418
rect 19378 23366 19390 23418
rect 19442 23366 28428 23418
rect 1104 23344 28428 23366
rect 3050 23304 3056 23316
rect 3011 23276 3056 23304
rect 3050 23264 3056 23276
rect 3108 23264 3114 23316
rect 5258 23264 5264 23316
rect 5316 23304 5322 23316
rect 9953 23307 10011 23313
rect 5316 23276 9628 23304
rect 5316 23264 5322 23276
rect 1854 23236 1860 23248
rect 1815 23208 1860 23236
rect 1854 23196 1860 23208
rect 1912 23196 1918 23248
rect 2777 23239 2835 23245
rect 2777 23205 2789 23239
rect 2823 23236 2835 23239
rect 3878 23236 3884 23248
rect 2823 23208 3884 23236
rect 2823 23205 2835 23208
rect 2777 23199 2835 23205
rect 3878 23196 3884 23208
rect 3936 23236 3942 23248
rect 9600 23236 9628 23276
rect 9953 23273 9965 23307
rect 9999 23304 10011 23307
rect 10410 23304 10416 23316
rect 9999 23276 10416 23304
rect 9999 23273 10011 23276
rect 9953 23267 10011 23273
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 10597 23307 10655 23313
rect 10597 23273 10609 23307
rect 10643 23304 10655 23307
rect 10962 23304 10968 23316
rect 10643 23276 10968 23304
rect 10643 23273 10655 23276
rect 10597 23267 10655 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 14921 23307 14979 23313
rect 14921 23273 14933 23307
rect 14967 23304 14979 23307
rect 15102 23304 15108 23316
rect 14967 23276 15108 23304
rect 14967 23273 14979 23276
rect 14921 23267 14979 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 16761 23307 16819 23313
rect 16761 23273 16773 23307
rect 16807 23304 16819 23307
rect 17310 23304 17316 23316
rect 16807 23276 17316 23304
rect 16807 23273 16819 23276
rect 16761 23267 16819 23273
rect 17310 23264 17316 23276
rect 17368 23264 17374 23316
rect 18414 23304 18420 23316
rect 18375 23276 18420 23304
rect 18414 23264 18420 23276
rect 18472 23264 18478 23316
rect 18690 23264 18696 23316
rect 18748 23304 18754 23316
rect 21174 23304 21180 23316
rect 18748 23276 21180 23304
rect 18748 23264 18754 23276
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 22738 23264 22744 23316
rect 22796 23304 22802 23316
rect 23477 23307 23535 23313
rect 23477 23304 23489 23307
rect 22796 23276 23489 23304
rect 22796 23264 22802 23276
rect 23477 23273 23489 23276
rect 23523 23273 23535 23307
rect 23477 23267 23535 23273
rect 26142 23264 26148 23316
rect 26200 23304 26206 23316
rect 27433 23307 27491 23313
rect 27433 23304 27445 23307
rect 26200 23276 27445 23304
rect 26200 23264 26206 23276
rect 27433 23273 27445 23276
rect 27479 23273 27491 23307
rect 27433 23267 27491 23273
rect 14458 23236 14464 23248
rect 3936 23208 9536 23236
rect 9600 23208 14464 23236
rect 3936 23196 3942 23208
rect 2498 23168 2504 23180
rect 2459 23140 2504 23168
rect 2498 23128 2504 23140
rect 2556 23128 2562 23180
rect 2590 23128 2596 23180
rect 2648 23168 2654 23180
rect 2685 23171 2743 23177
rect 2685 23168 2697 23171
rect 2648 23140 2697 23168
rect 2648 23128 2654 23140
rect 2685 23137 2697 23140
rect 2731 23137 2743 23171
rect 2685 23131 2743 23137
rect 2869 23171 2927 23177
rect 2869 23137 2881 23171
rect 2915 23168 2927 23171
rect 3142 23168 3148 23180
rect 2915 23140 3148 23168
rect 2915 23137 2927 23140
rect 2869 23131 2927 23137
rect 3142 23128 3148 23140
rect 3200 23128 3206 23180
rect 6638 23168 6644 23180
rect 6599 23140 6644 23168
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 9508 23177 9536 23208
rect 14458 23196 14464 23208
rect 14516 23196 14522 23248
rect 18137 23239 18195 23245
rect 18137 23236 18149 23239
rect 17972 23208 18149 23236
rect 8389 23171 8447 23177
rect 8389 23137 8401 23171
rect 8435 23137 8447 23171
rect 8389 23131 8447 23137
rect 9493 23171 9551 23177
rect 9493 23137 9505 23171
rect 9539 23137 9551 23171
rect 9493 23131 9551 23137
rect 5994 22992 6000 23044
rect 6052 23032 6058 23044
rect 7101 23035 7159 23041
rect 7101 23032 7113 23035
rect 6052 23004 7113 23032
rect 6052 22992 6058 23004
rect 7101 23001 7113 23004
rect 7147 23001 7159 23035
rect 8404 23032 8432 23131
rect 9674 23128 9680 23180
rect 9732 23168 9738 23180
rect 10505 23171 10563 23177
rect 10505 23168 10517 23171
rect 9732 23140 10517 23168
rect 9732 23128 9738 23140
rect 10505 23137 10517 23140
rect 10551 23137 10563 23171
rect 10505 23131 10563 23137
rect 11416 23171 11474 23177
rect 11416 23137 11428 23171
rect 11462 23168 11474 23171
rect 11974 23168 11980 23180
rect 11462 23140 11980 23168
rect 11462 23137 11474 23140
rect 11416 23131 11474 23137
rect 11974 23128 11980 23140
rect 12032 23128 12038 23180
rect 12986 23168 12992 23180
rect 12947 23140 12992 23168
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 13078 23128 13084 23180
rect 13136 23168 13142 23180
rect 13173 23171 13231 23177
rect 13173 23168 13185 23171
rect 13136 23140 13185 23168
rect 13136 23128 13142 23140
rect 13173 23137 13185 23140
rect 13219 23137 13231 23171
rect 13446 23168 13452 23180
rect 13407 23140 13452 23168
rect 13173 23131 13231 23137
rect 13446 23128 13452 23140
rect 13504 23128 13510 23180
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23168 13783 23171
rect 14182 23168 14188 23180
rect 13771 23140 14188 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 14826 23168 14832 23180
rect 14787 23140 14832 23168
rect 14826 23128 14832 23140
rect 14884 23128 14890 23180
rect 15654 23128 15660 23180
rect 15712 23168 15718 23180
rect 16025 23171 16083 23177
rect 16025 23168 16037 23171
rect 15712 23140 16037 23168
rect 15712 23128 15718 23140
rect 16025 23137 16037 23140
rect 16071 23137 16083 23171
rect 16206 23168 16212 23180
rect 16167 23140 16212 23168
rect 16025 23131 16083 23137
rect 16206 23128 16212 23140
rect 16264 23128 16270 23180
rect 16574 23168 16580 23180
rect 16535 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 17405 23171 17463 23177
rect 17405 23137 17417 23171
rect 17451 23137 17463 23171
rect 17862 23168 17868 23180
rect 17823 23140 17868 23168
rect 17405 23131 17463 23137
rect 10962 23060 10968 23112
rect 11020 23100 11026 23112
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 11020 23072 11161 23100
rect 11020 23060 11026 23072
rect 11149 23069 11161 23072
rect 11195 23069 11207 23103
rect 11149 23063 11207 23069
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 16301 23103 16359 23109
rect 16301 23100 16313 23103
rect 15068 23072 16313 23100
rect 15068 23060 15074 23072
rect 16301 23069 16313 23072
rect 16347 23069 16359 23103
rect 16301 23063 16359 23069
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23069 16451 23103
rect 16393 23063 16451 23069
rect 11054 23032 11060 23044
rect 8404 23004 11060 23032
rect 7101 22995 7159 23001
rect 11054 22992 11060 23004
rect 11112 22992 11118 23044
rect 13538 23032 13544 23044
rect 13499 23004 13544 23032
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 16022 22992 16028 23044
rect 16080 23032 16086 23044
rect 16408 23032 16436 23063
rect 17218 23032 17224 23044
rect 16080 23004 16436 23032
rect 17179 23004 17224 23032
rect 16080 22992 16086 23004
rect 17218 22992 17224 23004
rect 17276 22992 17282 23044
rect 1946 22964 1952 22976
rect 1907 22936 1952 22964
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 6825 22967 6883 22973
rect 6825 22933 6837 22967
rect 6871 22964 6883 22967
rect 6914 22964 6920 22976
rect 6871 22936 6920 22964
rect 6871 22933 6883 22936
rect 6825 22927 6883 22933
rect 6914 22924 6920 22936
rect 6972 22964 6978 22976
rect 8202 22964 8208 22976
rect 6972 22936 8208 22964
rect 6972 22924 6978 22936
rect 8202 22924 8208 22936
rect 8260 22964 8266 22976
rect 8573 22967 8631 22973
rect 8573 22964 8585 22967
rect 8260 22936 8585 22964
rect 8260 22924 8266 22936
rect 8573 22933 8585 22936
rect 8619 22964 8631 22967
rect 9585 22967 9643 22973
rect 9585 22964 9597 22967
rect 8619 22936 9597 22964
rect 8619 22933 8631 22936
rect 8573 22927 8631 22933
rect 9585 22933 9597 22936
rect 9631 22933 9643 22967
rect 9585 22927 9643 22933
rect 10502 22924 10508 22976
rect 10560 22964 10566 22976
rect 10870 22964 10876 22976
rect 10560 22936 10876 22964
rect 10560 22924 10566 22936
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 12066 22924 12072 22976
rect 12124 22964 12130 22976
rect 12529 22967 12587 22973
rect 12529 22964 12541 22967
rect 12124 22936 12541 22964
rect 12124 22924 12130 22936
rect 12529 22933 12541 22936
rect 12575 22933 12587 22967
rect 17420 22964 17448 23131
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 17972 23032 18000 23208
rect 18137 23205 18149 23208
rect 18183 23205 18195 23239
rect 18137 23199 18195 23205
rect 18782 23196 18788 23248
rect 18840 23236 18846 23248
rect 24302 23236 24308 23248
rect 18840 23208 24308 23236
rect 18840 23196 18846 23208
rect 24302 23196 24308 23208
rect 24360 23196 24366 23248
rect 26320 23239 26378 23245
rect 26320 23205 26332 23239
rect 26366 23236 26378 23239
rect 26694 23236 26700 23248
rect 26366 23208 26700 23236
rect 26366 23205 26378 23208
rect 26320 23199 26378 23205
rect 26694 23196 26700 23208
rect 26752 23196 26758 23248
rect 18049 23171 18107 23177
rect 18049 23137 18061 23171
rect 18095 23137 18107 23171
rect 18049 23131 18107 23137
rect 18064 23100 18092 23131
rect 18230 23128 18236 23180
rect 18288 23168 18294 23180
rect 18288 23140 18333 23168
rect 18288 23128 18294 23140
rect 18874 23128 18880 23180
rect 18932 23168 18938 23180
rect 19061 23171 19119 23177
rect 19061 23168 19073 23171
rect 18932 23140 19073 23168
rect 18932 23128 18938 23140
rect 19061 23137 19073 23140
rect 19107 23137 19119 23171
rect 20070 23168 20076 23180
rect 20031 23140 20076 23168
rect 19061 23131 19119 23137
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 20257 23171 20315 23177
rect 20257 23137 20269 23171
rect 20303 23137 20315 23171
rect 20257 23131 20315 23137
rect 20349 23171 20407 23177
rect 20349 23137 20361 23171
rect 20395 23137 20407 23171
rect 20349 23131 20407 23137
rect 18690 23100 18696 23112
rect 18064 23072 18696 23100
rect 18690 23060 18696 23072
rect 18748 23100 18754 23112
rect 20272 23100 20300 23131
rect 18748 23072 20300 23100
rect 20364 23100 20392 23131
rect 20438 23128 20444 23180
rect 20496 23168 20502 23180
rect 20496 23140 20541 23168
rect 20496 23128 20502 23140
rect 21634 23128 21640 23180
rect 21692 23168 21698 23180
rect 21801 23171 21859 23177
rect 21801 23168 21813 23171
rect 21692 23140 21813 23168
rect 21692 23128 21698 23140
rect 21801 23137 21813 23140
rect 21847 23137 21859 23171
rect 23385 23171 23443 23177
rect 23385 23168 23397 23171
rect 21801 23131 21859 23137
rect 22940 23140 23397 23168
rect 21450 23100 21456 23112
rect 20364 23072 21456 23100
rect 18748 23060 18754 23072
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 21542 23060 21548 23112
rect 21600 23100 21606 23112
rect 21600 23072 21645 23100
rect 21600 23060 21606 23072
rect 18138 23032 18144 23044
rect 17972 23004 18144 23032
rect 18138 22992 18144 23004
rect 18196 23032 18202 23044
rect 19518 23032 19524 23044
rect 18196 23004 19524 23032
rect 18196 22992 18202 23004
rect 19518 22992 19524 23004
rect 19576 22992 19582 23044
rect 20622 23032 20628 23044
rect 20583 23004 20628 23032
rect 20622 22992 20628 23004
rect 20680 22992 20686 23044
rect 18874 22964 18880 22976
rect 17420 22936 18880 22964
rect 12529 22927 12587 22933
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 21358 22924 21364 22976
rect 21416 22964 21422 22976
rect 22940 22973 22968 23140
rect 23385 23137 23397 23140
rect 23431 23137 23443 23171
rect 23385 23131 23443 23137
rect 24118 23128 24124 23180
rect 24176 23168 24182 23180
rect 24213 23171 24271 23177
rect 24213 23168 24225 23171
rect 24176 23140 24225 23168
rect 24176 23128 24182 23140
rect 24213 23137 24225 23140
rect 24259 23137 24271 23171
rect 24213 23131 24271 23137
rect 26050 23100 26056 23112
rect 24044 23072 26056 23100
rect 23474 22992 23480 23044
rect 23532 23032 23538 23044
rect 23934 23032 23940 23044
rect 23532 23004 23940 23032
rect 23532 22992 23538 23004
rect 23934 22992 23940 23004
rect 23992 23032 23998 23044
rect 24044 23041 24072 23072
rect 26050 23060 26056 23072
rect 26108 23060 26114 23112
rect 24029 23035 24087 23041
rect 24029 23032 24041 23035
rect 23992 23004 24041 23032
rect 23992 22992 23998 23004
rect 24029 23001 24041 23004
rect 24075 23001 24087 23035
rect 24029 22995 24087 23001
rect 22925 22967 22983 22973
rect 22925 22964 22937 22967
rect 21416 22936 22937 22964
rect 21416 22924 21422 22936
rect 22925 22933 22937 22936
rect 22971 22933 22983 22967
rect 22925 22927 22983 22933
rect 24302 22924 24308 22976
rect 24360 22964 24366 22976
rect 25314 22964 25320 22976
rect 24360 22936 25320 22964
rect 24360 22924 24366 22936
rect 25314 22924 25320 22936
rect 25372 22924 25378 22976
rect 1104 22874 28428 22896
rect 1104 22822 5536 22874
rect 5588 22822 5600 22874
rect 5652 22822 5664 22874
rect 5716 22822 5728 22874
rect 5780 22822 14644 22874
rect 14696 22822 14708 22874
rect 14760 22822 14772 22874
rect 14824 22822 14836 22874
rect 14888 22822 23752 22874
rect 23804 22822 23816 22874
rect 23868 22822 23880 22874
rect 23932 22822 23944 22874
rect 23996 22822 28428 22874
rect 1104 22800 28428 22822
rect 5166 22720 5172 22772
rect 5224 22760 5230 22772
rect 5721 22763 5779 22769
rect 5721 22760 5733 22763
rect 5224 22732 5733 22760
rect 5224 22720 5230 22732
rect 5721 22729 5733 22732
rect 5767 22729 5779 22763
rect 10410 22760 10416 22772
rect 10371 22732 10416 22760
rect 5721 22723 5779 22729
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 10594 22720 10600 22772
rect 10652 22760 10658 22772
rect 12161 22763 12219 22769
rect 12161 22760 12173 22763
rect 10652 22732 12173 22760
rect 10652 22720 10658 22732
rect 12161 22729 12173 22732
rect 12207 22729 12219 22763
rect 12161 22723 12219 22729
rect 14090 22720 14096 22772
rect 14148 22760 14154 22772
rect 14185 22763 14243 22769
rect 14185 22760 14197 22763
rect 14148 22732 14197 22760
rect 14148 22720 14154 22732
rect 14185 22729 14197 22732
rect 14231 22729 14243 22763
rect 14185 22723 14243 22729
rect 14829 22763 14887 22769
rect 14829 22729 14841 22763
rect 14875 22760 14887 22763
rect 15010 22760 15016 22772
rect 14875 22732 15016 22760
rect 14875 22729 14887 22732
rect 14829 22723 14887 22729
rect 1946 22652 1952 22704
rect 2004 22692 2010 22704
rect 2004 22664 11008 22692
rect 2004 22652 2010 22664
rect 7374 22624 7380 22636
rect 7208 22596 7380 22624
rect 1857 22559 1915 22565
rect 1857 22525 1869 22559
rect 1903 22556 1915 22559
rect 5258 22556 5264 22568
rect 1903 22528 5264 22556
rect 1903 22525 1915 22528
rect 1857 22519 1915 22525
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 5905 22559 5963 22565
rect 5905 22525 5917 22559
rect 5951 22556 5963 22559
rect 6270 22556 6276 22568
rect 5951 22528 6276 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 6270 22516 6276 22528
rect 6328 22516 6334 22568
rect 6822 22556 6828 22568
rect 6783 22528 6828 22556
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 7208 22565 7236 22596
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 10980 22624 11008 22664
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 11112 22664 12434 22692
rect 11112 22652 11118 22664
rect 12250 22624 12256 22636
rect 9732 22596 10364 22624
rect 10980 22596 12256 22624
rect 9732 22584 9738 22596
rect 7009 22559 7067 22565
rect 7009 22525 7021 22559
rect 7055 22525 7067 22559
rect 7009 22519 7067 22525
rect 7193 22559 7251 22565
rect 7193 22525 7205 22559
rect 7239 22525 7251 22559
rect 7193 22519 7251 22525
rect 2038 22488 2044 22500
rect 1999 22460 2044 22488
rect 2038 22448 2044 22460
rect 2096 22448 2102 22500
rect 7024 22432 7052 22519
rect 7282 22516 7288 22568
rect 7340 22556 7346 22568
rect 7558 22556 7564 22568
rect 7340 22528 7564 22556
rect 7340 22516 7346 22528
rect 7558 22516 7564 22528
rect 7616 22556 7622 22568
rect 7837 22559 7895 22565
rect 7837 22556 7849 22559
rect 7616 22528 7849 22556
rect 7616 22516 7622 22528
rect 7837 22525 7849 22528
rect 7883 22525 7895 22559
rect 8938 22556 8944 22568
rect 8899 22528 8944 22556
rect 7837 22519 7895 22525
rect 8938 22516 8944 22528
rect 8996 22516 9002 22568
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 10060 22565 10088 22596
rect 9861 22559 9919 22565
rect 9861 22556 9873 22559
rect 9180 22528 9873 22556
rect 9180 22516 9186 22528
rect 9861 22525 9873 22528
rect 9907 22525 9919 22559
rect 9861 22519 9919 22525
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22525 10103 22559
rect 10226 22556 10232 22568
rect 10187 22528 10232 22556
rect 10045 22519 10103 22525
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 10336 22556 10364 22596
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 12406 22624 12434 22664
rect 13814 22652 13820 22704
rect 13872 22692 13878 22704
rect 14844 22692 14872 22723
rect 15010 22720 15016 22732
rect 15068 22720 15074 22772
rect 26789 22763 26847 22769
rect 26789 22760 26801 22763
rect 15120 22732 26801 22760
rect 13872 22664 14872 22692
rect 13872 22652 13878 22664
rect 12406 22596 12940 22624
rect 11057 22559 11115 22565
rect 10336 22528 11008 22556
rect 7098 22448 7104 22500
rect 7156 22488 7162 22500
rect 9582 22488 9588 22500
rect 7156 22460 7201 22488
rect 7254 22460 9588 22488
rect 7156 22448 7162 22460
rect 7006 22380 7012 22432
rect 7064 22420 7070 22432
rect 7254 22420 7282 22460
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 10137 22491 10195 22497
rect 10137 22457 10149 22491
rect 10183 22457 10195 22491
rect 10594 22488 10600 22500
rect 10137 22451 10195 22457
rect 10336 22460 10600 22488
rect 7374 22420 7380 22432
rect 7064 22392 7282 22420
rect 7335 22392 7380 22420
rect 7064 22380 7070 22392
rect 7374 22380 7380 22392
rect 7432 22380 7438 22432
rect 7929 22423 7987 22429
rect 7929 22389 7941 22423
rect 7975 22420 7987 22423
rect 8846 22420 8852 22432
rect 7975 22392 8852 22420
rect 7975 22389 7987 22392
rect 7929 22383 7987 22389
rect 8846 22380 8852 22392
rect 8904 22380 8910 22432
rect 9033 22423 9091 22429
rect 9033 22389 9045 22423
rect 9079 22420 9091 22423
rect 9214 22420 9220 22432
rect 9079 22392 9220 22420
rect 9079 22389 9091 22392
rect 9033 22383 9091 22389
rect 9214 22380 9220 22392
rect 9272 22380 9278 22432
rect 10152 22420 10180 22451
rect 10336 22420 10364 22460
rect 10594 22448 10600 22460
rect 10652 22448 10658 22500
rect 10980 22488 11008 22528
rect 11057 22525 11069 22559
rect 11103 22556 11115 22559
rect 11606 22556 11612 22568
rect 11103 22528 11612 22556
rect 11103 22525 11115 22528
rect 11057 22519 11115 22525
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 12066 22556 12072 22568
rect 12027 22528 12072 22556
rect 12066 22516 12072 22528
rect 12124 22516 12130 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 12805 22559 12863 22565
rect 12805 22556 12817 22559
rect 12768 22528 12817 22556
rect 12768 22516 12774 22528
rect 12805 22525 12817 22528
rect 12851 22525 12863 22559
rect 12912 22556 12940 22596
rect 14645 22559 14703 22565
rect 14645 22556 14657 22559
rect 12912 22528 14657 22556
rect 12805 22519 12863 22525
rect 14645 22525 14657 22528
rect 14691 22525 14703 22559
rect 14645 22519 14703 22525
rect 13072 22491 13130 22497
rect 10980 22460 13032 22488
rect 10152 22392 10364 22420
rect 10873 22423 10931 22429
rect 10873 22389 10885 22423
rect 10919 22420 10931 22423
rect 11146 22420 11152 22432
rect 10919 22392 11152 22420
rect 10919 22389 10931 22392
rect 10873 22383 10931 22389
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 13004 22420 13032 22460
rect 13072 22457 13084 22491
rect 13118 22488 13130 22491
rect 13630 22488 13636 22500
rect 13118 22460 13636 22488
rect 13118 22457 13130 22460
rect 13072 22451 13130 22457
rect 13630 22448 13636 22460
rect 13688 22448 13694 22500
rect 15120 22420 15148 22732
rect 26789 22729 26801 22732
rect 26835 22729 26847 22763
rect 26789 22723 26847 22729
rect 15470 22652 15476 22704
rect 15528 22692 15534 22704
rect 15657 22695 15715 22701
rect 15657 22692 15669 22695
rect 15528 22664 15669 22692
rect 15528 22652 15534 22664
rect 15657 22661 15669 22664
rect 15703 22661 15715 22695
rect 16390 22692 16396 22704
rect 16351 22664 16396 22692
rect 15657 22655 15715 22661
rect 16390 22652 16396 22664
rect 16448 22652 16454 22704
rect 21637 22695 21695 22701
rect 17144 22664 18000 22692
rect 15470 22516 15476 22568
rect 15528 22556 15534 22568
rect 17144 22556 17172 22664
rect 17862 22624 17868 22636
rect 17328 22596 17868 22624
rect 17328 22568 17356 22596
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 17972 22624 18000 22664
rect 21637 22661 21649 22695
rect 21683 22661 21695 22695
rect 21637 22655 21695 22661
rect 20530 22624 20536 22636
rect 17972 22596 18828 22624
rect 17310 22556 17316 22568
rect 15528 22528 17172 22556
rect 17223 22528 17316 22556
rect 15528 22516 15534 22528
rect 17310 22516 17316 22528
rect 17368 22516 17374 22568
rect 17586 22556 17592 22568
rect 17547 22528 17592 22556
rect 17586 22516 17592 22528
rect 17644 22516 17650 22568
rect 17678 22516 17684 22568
rect 17736 22556 17742 22568
rect 18230 22556 18236 22568
rect 17736 22528 18236 22556
rect 17736 22516 17742 22528
rect 18230 22516 18236 22528
rect 18288 22516 18294 22568
rect 18322 22516 18328 22568
rect 18380 22556 18386 22568
rect 18693 22559 18751 22565
rect 18693 22556 18705 22559
rect 18380 22528 18705 22556
rect 18380 22516 18386 22528
rect 18693 22525 18705 22528
rect 18739 22525 18751 22559
rect 18800 22556 18828 22596
rect 19996 22596 20536 22624
rect 19996 22556 20024 22596
rect 20530 22584 20536 22596
rect 20588 22584 20594 22636
rect 21652 22568 21680 22655
rect 22186 22652 22192 22704
rect 22244 22692 22250 22704
rect 23290 22692 23296 22704
rect 22244 22664 23296 22692
rect 22244 22652 22250 22664
rect 23290 22652 23296 22664
rect 23348 22692 23354 22704
rect 23934 22692 23940 22704
rect 23348 22664 23940 22692
rect 23348 22652 23354 22664
rect 23934 22652 23940 22664
rect 23992 22652 23998 22704
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 21968 22596 22968 22624
rect 21968 22584 21974 22596
rect 18800 22528 20024 22556
rect 18693 22519 18751 22525
rect 20070 22516 20076 22568
rect 20128 22556 20134 22568
rect 21085 22559 21143 22565
rect 21085 22556 21097 22559
rect 20128 22528 21097 22556
rect 20128 22516 20134 22528
rect 21085 22525 21097 22528
rect 21131 22525 21143 22559
rect 21358 22556 21364 22568
rect 21319 22528 21364 22556
rect 21085 22519 21143 22525
rect 16114 22448 16120 22500
rect 16172 22488 16178 22500
rect 16209 22491 16267 22497
rect 16209 22488 16221 22491
rect 16172 22460 16221 22488
rect 16172 22448 16178 22460
rect 16209 22457 16221 22460
rect 16255 22457 16267 22491
rect 16209 22451 16267 22457
rect 17402 22448 17408 22500
rect 17460 22488 17466 22500
rect 17497 22491 17555 22497
rect 17497 22488 17509 22491
rect 17460 22460 17509 22488
rect 17460 22448 17466 22460
rect 17497 22457 17509 22460
rect 17543 22457 17555 22491
rect 17497 22451 17555 22457
rect 18414 22448 18420 22500
rect 18472 22488 18478 22500
rect 18938 22491 18996 22497
rect 18938 22488 18950 22491
rect 18472 22460 18950 22488
rect 18472 22448 18478 22460
rect 18938 22457 18950 22460
rect 18984 22457 18996 22491
rect 18938 22451 18996 22457
rect 19150 22448 19156 22500
rect 19208 22488 19214 22500
rect 19978 22488 19984 22500
rect 19208 22460 19984 22488
rect 19208 22448 19214 22460
rect 19978 22448 19984 22460
rect 20036 22448 20042 22500
rect 17862 22420 17868 22432
rect 13004 22392 15148 22420
rect 17823 22392 17868 22420
rect 17862 22380 17868 22392
rect 17920 22380 17926 22432
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18782 22420 18788 22432
rect 18104 22392 18788 22420
rect 18104 22380 18110 22392
rect 18782 22380 18788 22392
rect 18840 22380 18846 22432
rect 19794 22380 19800 22432
rect 19852 22420 19858 22432
rect 20073 22423 20131 22429
rect 20073 22420 20085 22423
rect 19852 22392 20085 22420
rect 19852 22380 19858 22392
rect 20073 22389 20085 22392
rect 20119 22420 20131 22423
rect 20622 22420 20628 22432
rect 20119 22392 20628 22420
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 21100 22420 21128 22519
rect 21358 22516 21364 22528
rect 21416 22516 21422 22568
rect 21450 22516 21456 22568
rect 21508 22565 21514 22568
rect 21508 22559 21535 22565
rect 21523 22525 21535 22559
rect 21508 22519 21535 22525
rect 21508 22516 21514 22519
rect 21634 22516 21640 22568
rect 21692 22516 21698 22568
rect 22940 22565 22968 22596
rect 23474 22584 23480 22636
rect 23532 22624 23538 22636
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23532 22596 24041 22624
rect 23532 22584 23538 22596
rect 24029 22593 24041 22596
rect 24075 22593 24087 22627
rect 26053 22627 26111 22633
rect 26053 22624 26065 22627
rect 24029 22587 24087 22593
rect 25332 22596 26065 22624
rect 22557 22559 22615 22565
rect 22557 22525 22569 22559
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 22925 22559 22983 22565
rect 22925 22525 22937 22559
rect 22971 22525 22983 22559
rect 22925 22519 22983 22525
rect 21266 22488 21272 22500
rect 21227 22460 21272 22488
rect 21266 22448 21272 22460
rect 21324 22448 21330 22500
rect 22572 22488 22600 22519
rect 24578 22516 24584 22568
rect 24636 22556 24642 22568
rect 25332 22556 25360 22596
rect 26053 22593 26065 22596
rect 26099 22593 26111 22627
rect 26053 22587 26111 22593
rect 24636 22528 25360 22556
rect 25961 22559 26019 22565
rect 24636 22516 24642 22528
rect 25961 22525 25973 22559
rect 26007 22556 26019 22559
rect 26142 22556 26148 22568
rect 26007 22528 26148 22556
rect 26007 22525 26019 22528
rect 25961 22519 26019 22525
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 26697 22559 26755 22565
rect 26697 22525 26709 22559
rect 26743 22556 26755 22559
rect 26786 22556 26792 22568
rect 26743 22528 26792 22556
rect 26743 22525 26755 22528
rect 26697 22519 26755 22525
rect 26786 22516 26792 22528
rect 26844 22516 26850 22568
rect 21816 22460 22600 22488
rect 21816 22420 21844 22460
rect 22646 22448 22652 22500
rect 22704 22488 22710 22500
rect 22741 22491 22799 22497
rect 22741 22488 22753 22491
rect 22704 22460 22753 22488
rect 22704 22448 22710 22460
rect 22741 22457 22753 22460
rect 22787 22457 22799 22491
rect 22741 22451 22799 22457
rect 22833 22491 22891 22497
rect 22833 22457 22845 22491
rect 22879 22488 22891 22491
rect 24296 22491 24354 22497
rect 22879 22460 22968 22488
rect 22879 22457 22891 22460
rect 22833 22451 22891 22457
rect 21100 22392 21844 22420
rect 22554 22380 22560 22432
rect 22612 22420 22618 22432
rect 22940 22420 22968 22460
rect 24296 22457 24308 22491
rect 24342 22488 24354 22491
rect 25774 22488 25780 22500
rect 24342 22460 25780 22488
rect 24342 22457 24354 22460
rect 24296 22451 24354 22457
rect 25774 22448 25780 22460
rect 25832 22448 25838 22500
rect 23106 22420 23112 22432
rect 22612 22392 22968 22420
rect 23067 22392 23112 22420
rect 22612 22380 22618 22392
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 25406 22420 25412 22432
rect 25367 22392 25412 22420
rect 25406 22380 25412 22392
rect 25464 22380 25470 22432
rect 1104 22330 28428 22352
rect 1104 22278 10090 22330
rect 10142 22278 10154 22330
rect 10206 22278 10218 22330
rect 10270 22278 10282 22330
rect 10334 22278 19198 22330
rect 19250 22278 19262 22330
rect 19314 22278 19326 22330
rect 19378 22278 19390 22330
rect 19442 22278 28428 22330
rect 1104 22256 28428 22278
rect 6638 22216 6644 22228
rect 5644 22188 6644 22216
rect 5166 22040 5172 22092
rect 5224 22080 5230 22092
rect 5644 22089 5672 22188
rect 6638 22176 6644 22188
rect 6696 22176 6702 22228
rect 6822 22176 6828 22228
rect 6880 22176 6886 22228
rect 6914 22176 6920 22228
rect 6972 22176 6978 22228
rect 7009 22219 7067 22225
rect 7009 22185 7021 22219
rect 7055 22216 7067 22219
rect 7282 22216 7288 22228
rect 7055 22188 7288 22216
rect 7055 22185 7067 22188
rect 7009 22179 7067 22185
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 11974 22216 11980 22228
rect 11935 22188 11980 22216
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12437 22219 12495 22225
rect 12437 22185 12449 22219
rect 12483 22216 12495 22219
rect 12710 22216 12716 22228
rect 12483 22188 12716 22216
rect 12483 22185 12495 22188
rect 12437 22179 12495 22185
rect 12710 22176 12716 22188
rect 12768 22176 12774 22228
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 17034 22216 17040 22228
rect 13504 22188 17040 22216
rect 13504 22176 13510 22188
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 17586 22216 17592 22228
rect 17547 22188 17592 22216
rect 17586 22176 17592 22188
rect 17644 22176 17650 22228
rect 18414 22176 18420 22228
rect 18472 22216 18478 22228
rect 19061 22219 19119 22225
rect 19061 22216 19073 22219
rect 18472 22188 19073 22216
rect 18472 22176 18478 22188
rect 19061 22185 19073 22188
rect 19107 22185 19119 22219
rect 19061 22179 19119 22185
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 22922 22216 22928 22228
rect 22704 22188 22928 22216
rect 22704 22176 22710 22188
rect 22922 22176 22928 22188
rect 22980 22216 22986 22228
rect 22980 22188 23704 22216
rect 22980 22176 22986 22188
rect 6454 22108 6460 22160
rect 6512 22148 6518 22160
rect 6840 22148 6868 22176
rect 6512 22120 6868 22148
rect 6932 22148 6960 22176
rect 7653 22151 7711 22157
rect 7653 22148 7665 22151
rect 6932 22120 7665 22148
rect 6512 22108 6518 22120
rect 6840 22094 6868 22120
rect 7653 22117 7665 22120
rect 7699 22148 7711 22151
rect 10686 22148 10692 22160
rect 7699 22120 8953 22148
rect 7699 22117 7711 22120
rect 7653 22111 7711 22117
rect 5629 22083 5687 22089
rect 5629 22080 5641 22083
rect 5224 22052 5641 22080
rect 5224 22040 5230 22052
rect 5629 22049 5641 22052
rect 5675 22049 5687 22083
rect 5629 22043 5687 22049
rect 5896 22083 5954 22089
rect 5896 22049 5908 22083
rect 5942 22080 5954 22083
rect 6840 22080 6914 22094
rect 7469 22083 7527 22089
rect 7469 22080 7481 22083
rect 5942 22052 6684 22080
rect 6840 22066 7481 22080
rect 6886 22052 7481 22066
rect 5942 22049 5954 22052
rect 5896 22043 5954 22049
rect 6656 21944 6684 22052
rect 7469 22049 7481 22052
rect 7515 22049 7527 22083
rect 7469 22043 7527 22049
rect 7558 22040 7564 22092
rect 7616 22080 7622 22092
rect 7745 22083 7803 22089
rect 7745 22080 7757 22083
rect 7616 22052 7757 22080
rect 7616 22040 7622 22052
rect 7745 22049 7757 22052
rect 7791 22049 7803 22083
rect 7745 22043 7803 22049
rect 7837 22083 7895 22089
rect 7837 22049 7849 22083
rect 7883 22049 7895 22083
rect 7837 22043 7895 22049
rect 6730 21972 6736 22024
rect 6788 22012 6794 22024
rect 7190 22012 7196 22024
rect 6788 21984 7196 22012
rect 6788 21972 6794 21984
rect 7190 21972 7196 21984
rect 7248 22012 7254 22024
rect 7852 22012 7880 22043
rect 7248 21984 7880 22012
rect 8925 22012 8953 22120
rect 9692 22120 10692 22148
rect 9122 22040 9128 22092
rect 9180 22080 9186 22092
rect 9493 22083 9551 22089
rect 9493 22080 9505 22083
rect 9180 22052 9505 22080
rect 9180 22040 9186 22052
rect 9493 22049 9505 22052
rect 9539 22049 9551 22083
rect 9493 22043 9551 22049
rect 9582 22040 9588 22092
rect 9640 22080 9646 22092
rect 9692 22089 9720 22120
rect 10686 22108 10692 22120
rect 10744 22108 10750 22160
rect 11701 22151 11759 22157
rect 11701 22117 11713 22151
rect 11747 22148 11759 22151
rect 12066 22148 12072 22160
rect 11747 22120 12072 22148
rect 11747 22117 11759 22120
rect 11701 22111 11759 22117
rect 12066 22108 12072 22120
rect 12124 22108 12130 22160
rect 15657 22151 15715 22157
rect 15657 22148 15669 22151
rect 12544 22120 15669 22148
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 9640 22052 9689 22080
rect 9640 22040 9646 22052
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 9765 22083 9823 22089
rect 9765 22049 9777 22083
rect 9811 22049 9823 22083
rect 9765 22043 9823 22049
rect 9861 22083 9919 22089
rect 9861 22049 9873 22083
rect 9907 22080 9919 22083
rect 10042 22080 10048 22092
rect 9907 22052 10048 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 8925 21984 9674 22012
rect 7248 21972 7254 21984
rect 9646 21956 9674 21984
rect 9775 21956 9803 22043
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 10505 22083 10563 22089
rect 10505 22049 10517 22083
rect 10551 22080 10563 22083
rect 10594 22080 10600 22092
rect 10551 22052 10600 22080
rect 10551 22049 10563 22052
rect 10505 22043 10563 22049
rect 10594 22040 10600 22052
rect 10652 22080 10658 22092
rect 10870 22080 10876 22092
rect 10652 22052 10876 22080
rect 10652 22040 10658 22052
rect 10870 22040 10876 22052
rect 10928 22040 10934 22092
rect 11422 22080 11428 22092
rect 11383 22052 11428 22080
rect 11422 22040 11428 22052
rect 11480 22040 11486 22092
rect 11609 22083 11667 22089
rect 11609 22049 11621 22083
rect 11655 22049 11667 22083
rect 11609 22043 11667 22049
rect 11793 22083 11851 22089
rect 11793 22049 11805 22083
rect 11839 22080 11851 22083
rect 12544 22080 12572 22120
rect 15657 22117 15669 22120
rect 15703 22148 15715 22151
rect 15930 22148 15936 22160
rect 15703 22120 15936 22148
rect 15703 22117 15715 22120
rect 15657 22111 15715 22117
rect 15930 22108 15936 22120
rect 15988 22108 15994 22160
rect 19242 22148 19248 22160
rect 18524 22120 19248 22148
rect 11839 22052 12572 22080
rect 12621 22083 12679 22089
rect 11839 22049 11851 22052
rect 11793 22043 11851 22049
rect 12621 22049 12633 22083
rect 12667 22049 12679 22083
rect 12621 22043 12679 22049
rect 8021 21947 8079 21953
rect 8021 21944 8033 21947
rect 6656 21916 8033 21944
rect 8021 21913 8033 21916
rect 8067 21913 8079 21947
rect 9646 21916 9680 21956
rect 8021 21907 8079 21913
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 9766 21904 9772 21956
rect 9824 21944 9830 21956
rect 10686 21944 10692 21956
rect 9824 21916 10692 21944
rect 9824 21904 9830 21916
rect 10686 21904 10692 21916
rect 10744 21904 10750 21956
rect 11624 21944 11652 22043
rect 11698 21972 11704 22024
rect 11756 22012 11762 22024
rect 12636 22012 12664 22043
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 13449 22083 13507 22089
rect 13449 22080 13461 22083
rect 13044 22052 13461 22080
rect 13044 22040 13050 22052
rect 13449 22049 13461 22052
rect 13495 22049 13507 22083
rect 13449 22043 13507 22049
rect 14737 22083 14795 22089
rect 14737 22049 14749 22083
rect 14783 22080 14795 22083
rect 15286 22080 15292 22092
rect 14783 22052 15292 22080
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 15286 22040 15292 22052
rect 15344 22040 15350 22092
rect 15473 22083 15531 22089
rect 15473 22049 15485 22083
rect 15519 22080 15531 22083
rect 15838 22080 15844 22092
rect 15519 22052 15844 22080
rect 15519 22049 15531 22052
rect 15473 22043 15531 22049
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 16476 22083 16534 22089
rect 16476 22049 16488 22083
rect 16522 22080 16534 22083
rect 17862 22080 17868 22092
rect 16522 22052 17868 22080
rect 16522 22049 16534 22052
rect 16476 22043 16534 22049
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18524 22089 18552 22120
rect 19242 22108 19248 22120
rect 19300 22108 19306 22160
rect 19904 22120 20484 22148
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22049 18567 22083
rect 18509 22043 18567 22049
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22049 18751 22083
rect 18693 22043 18751 22049
rect 18785 22083 18843 22089
rect 18785 22049 18797 22083
rect 18831 22049 18843 22083
rect 18785 22043 18843 22049
rect 18877 22083 18935 22089
rect 18877 22049 18889 22083
rect 18923 22080 18935 22083
rect 19904 22080 19932 22120
rect 20456 22092 20484 22120
rect 20530 22108 20536 22160
rect 20588 22148 20594 22160
rect 21085 22151 21143 22157
rect 21085 22148 21097 22151
rect 20588 22120 21097 22148
rect 20588 22108 20594 22120
rect 21085 22117 21097 22120
rect 21131 22117 21143 22151
rect 21085 22111 21143 22117
rect 21269 22151 21327 22157
rect 21269 22117 21281 22151
rect 21315 22148 21327 22151
rect 21450 22148 21456 22160
rect 21315 22120 21456 22148
rect 21315 22117 21327 22120
rect 21269 22111 21327 22117
rect 18923 22052 19932 22080
rect 19981 22083 20039 22089
rect 18923 22049 18935 22052
rect 18877 22043 18935 22049
rect 19981 22049 19993 22083
rect 20027 22049 20039 22083
rect 19981 22043 20039 22049
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22049 20223 22083
rect 20165 22043 20223 22049
rect 16206 22012 16212 22024
rect 11756 21984 12664 22012
rect 16167 21984 16212 22012
rect 11756 21972 11762 21984
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 17402 21972 17408 22024
rect 17460 22012 17466 22024
rect 18708 22012 18736 22043
rect 17460 21984 18736 22012
rect 18800 22012 18828 22043
rect 19794 22012 19800 22024
rect 18800 21984 19800 22012
rect 17460 21972 17466 21984
rect 19794 21972 19800 21984
rect 19852 21972 19858 22024
rect 13262 21944 13268 21956
rect 11624 21916 13268 21944
rect 13262 21904 13268 21916
rect 13320 21904 13326 21956
rect 18322 21904 18328 21956
rect 18380 21944 18386 21956
rect 18966 21944 18972 21956
rect 18380 21916 18972 21944
rect 18380 21904 18386 21916
rect 18966 21904 18972 21916
rect 19024 21904 19030 21956
rect 19242 21904 19248 21956
rect 19300 21944 19306 21956
rect 19996 21944 20024 22043
rect 20180 21956 20208 22043
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 20438 22089 20444 22092
rect 20395 22083 20444 22089
rect 20312 22052 20357 22080
rect 20312 22040 20318 22052
rect 20395 22049 20407 22083
rect 20441 22049 20444 22083
rect 20395 22043 20444 22049
rect 20438 22040 20444 22043
rect 20496 22080 20502 22092
rect 21284 22080 21312 22111
rect 21450 22108 21456 22120
rect 21508 22148 21514 22160
rect 21910 22148 21916 22160
rect 21508 22120 21916 22148
rect 21508 22108 21514 22120
rect 21910 22108 21916 22120
rect 21968 22108 21974 22160
rect 22088 22151 22146 22157
rect 22088 22117 22100 22151
rect 22134 22148 22146 22151
rect 23106 22148 23112 22160
rect 22134 22120 23112 22148
rect 22134 22117 22146 22120
rect 22088 22111 22146 22117
rect 23106 22108 23112 22120
rect 23164 22108 23170 22160
rect 23676 22148 23704 22188
rect 24394 22176 24400 22228
rect 24452 22216 24458 22228
rect 25406 22216 25412 22228
rect 24452 22188 25412 22216
rect 24452 22176 24458 22188
rect 25406 22176 25412 22188
rect 25464 22216 25470 22228
rect 25774 22216 25780 22228
rect 25464 22188 25544 22216
rect 25735 22188 25780 22216
rect 25464 22176 25470 22188
rect 25516 22157 25544 22188
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 25501 22151 25559 22157
rect 23676 22120 25452 22148
rect 20496 22052 21312 22080
rect 20496 22040 20502 22052
rect 21542 22040 21548 22092
rect 21600 22080 21606 22092
rect 21821 22083 21879 22089
rect 21821 22080 21833 22083
rect 21600 22052 21833 22080
rect 21600 22040 21606 22052
rect 21821 22049 21833 22052
rect 21867 22080 21879 22083
rect 23474 22080 23480 22092
rect 21867 22052 23480 22080
rect 21867 22049 21879 22052
rect 21821 22043 21879 22049
rect 23474 22040 23480 22052
rect 23532 22040 23538 22092
rect 23566 22040 23572 22092
rect 23624 22080 23630 22092
rect 23661 22083 23719 22089
rect 23661 22080 23673 22083
rect 23624 22052 23673 22080
rect 23624 22040 23630 22052
rect 23661 22049 23673 22052
rect 23707 22049 23719 22083
rect 23842 22080 23848 22092
rect 23803 22052 23848 22080
rect 23661 22043 23719 22049
rect 23842 22040 23848 22052
rect 23900 22040 23906 22092
rect 23934 22040 23940 22092
rect 23992 22080 23998 22092
rect 24213 22083 24271 22089
rect 23992 22052 24037 22080
rect 23992 22040 23998 22052
rect 24213 22049 24225 22083
rect 24259 22080 24271 22083
rect 24762 22080 24768 22092
rect 24259 22052 24768 22080
rect 24259 22049 24271 22052
rect 24213 22043 24271 22049
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 25222 22080 25228 22092
rect 25183 22052 25228 22080
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 25424 22089 25452 22120
rect 25501 22117 25513 22151
rect 25547 22117 25559 22151
rect 25501 22111 25559 22117
rect 26789 22151 26847 22157
rect 26789 22117 26801 22151
rect 26835 22148 26847 22151
rect 27246 22148 27252 22160
rect 26835 22120 27252 22148
rect 26835 22117 26847 22120
rect 26789 22111 26847 22117
rect 27246 22108 27252 22120
rect 27304 22108 27310 22160
rect 27522 22148 27528 22160
rect 27483 22120 27528 22148
rect 27522 22108 27528 22120
rect 27580 22108 27586 22160
rect 25409 22083 25467 22089
rect 25409 22049 25421 22083
rect 25455 22049 25467 22083
rect 25409 22043 25467 22049
rect 25593 22083 25651 22089
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 25682 22080 25688 22092
rect 25639 22052 25688 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 26970 22080 26976 22092
rect 26931 22052 26976 22080
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 20070 21944 20076 21956
rect 19300 21916 20076 21944
rect 19300 21904 19306 21916
rect 20070 21904 20076 21916
rect 20128 21904 20134 21956
rect 20162 21904 20168 21956
rect 20220 21904 20226 21956
rect 23382 21904 23388 21956
rect 23440 21944 23446 21956
rect 23440 21916 23796 21944
rect 23440 21904 23446 21916
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 6730 21876 6736 21888
rect 6604 21848 6736 21876
rect 6604 21836 6610 21848
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 7190 21836 7196 21888
rect 7248 21876 7254 21888
rect 8110 21876 8116 21888
rect 7248 21848 8116 21876
rect 7248 21836 7254 21848
rect 8110 21836 8116 21848
rect 8168 21836 8174 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 10045 21879 10103 21885
rect 10045 21876 10057 21879
rect 10008 21848 10057 21876
rect 10008 21836 10014 21848
rect 10045 21845 10057 21848
rect 10091 21845 10103 21879
rect 10045 21839 10103 21845
rect 10502 21836 10508 21888
rect 10560 21876 10566 21888
rect 10597 21879 10655 21885
rect 10597 21876 10609 21879
rect 10560 21848 10609 21876
rect 10560 21836 10566 21848
rect 10597 21845 10609 21848
rect 10643 21845 10655 21879
rect 10597 21839 10655 21845
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 11698 21876 11704 21888
rect 11204 21848 11704 21876
rect 11204 21836 11210 21848
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 12802 21836 12808 21888
rect 12860 21876 12866 21888
rect 12986 21876 12992 21888
rect 12860 21848 12992 21876
rect 12860 21836 12866 21848
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 13541 21879 13599 21885
rect 13541 21876 13553 21879
rect 13504 21848 13553 21876
rect 13504 21836 13510 21848
rect 13541 21845 13553 21848
rect 13587 21845 13599 21879
rect 13541 21839 13599 21845
rect 13722 21836 13728 21888
rect 13780 21876 13786 21888
rect 14829 21879 14887 21885
rect 14829 21876 14841 21879
rect 13780 21848 14841 21876
rect 13780 21836 13786 21848
rect 14829 21845 14841 21848
rect 14875 21876 14887 21879
rect 15194 21876 15200 21888
rect 14875 21848 15200 21876
rect 14875 21845 14887 21848
rect 14829 21839 14887 21845
rect 15194 21836 15200 21848
rect 15252 21836 15258 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 15470 21876 15476 21888
rect 15344 21848 15476 21876
rect 15344 21836 15350 21848
rect 15470 21836 15476 21848
rect 15528 21836 15534 21888
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 18690 21876 18696 21888
rect 17368 21848 18696 21876
rect 17368 21836 17374 21848
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 20530 21876 20536 21888
rect 20491 21848 20536 21876
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 23201 21879 23259 21885
rect 23201 21876 23213 21879
rect 22612 21848 23213 21876
rect 22612 21836 22618 21848
rect 23201 21845 23213 21848
rect 23247 21845 23259 21879
rect 23201 21839 23259 21845
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 23661 21879 23719 21885
rect 23661 21876 23673 21879
rect 23624 21848 23673 21876
rect 23624 21836 23630 21848
rect 23661 21845 23673 21848
rect 23707 21845 23719 21879
rect 23768 21876 23796 21916
rect 23842 21904 23848 21956
rect 23900 21944 23906 21956
rect 25406 21944 25412 21956
rect 23900 21916 25412 21944
rect 23900 21904 23906 21916
rect 25406 21904 25412 21916
rect 25464 21904 25470 21956
rect 24121 21879 24179 21885
rect 24121 21876 24133 21879
rect 23768 21848 24133 21876
rect 23661 21839 23719 21845
rect 24121 21845 24133 21848
rect 24167 21845 24179 21879
rect 27614 21876 27620 21888
rect 27575 21848 27620 21876
rect 24121 21839 24179 21845
rect 27614 21836 27620 21848
rect 27672 21836 27678 21888
rect 1104 21786 28428 21808
rect 1104 21734 5536 21786
rect 5588 21734 5600 21786
rect 5652 21734 5664 21786
rect 5716 21734 5728 21786
rect 5780 21734 14644 21786
rect 14696 21734 14708 21786
rect 14760 21734 14772 21786
rect 14824 21734 14836 21786
rect 14888 21734 23752 21786
rect 23804 21734 23816 21786
rect 23868 21734 23880 21786
rect 23932 21734 23944 21786
rect 23996 21734 28428 21786
rect 1104 21712 28428 21734
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 6730 21672 6736 21684
rect 2271 21644 6736 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 6730 21632 6736 21644
rect 6788 21632 6794 21684
rect 7098 21632 7104 21684
rect 7156 21672 7162 21684
rect 8202 21672 8208 21684
rect 7156 21644 8208 21672
rect 7156 21632 7162 21644
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 8536 21644 10640 21672
rect 8536 21632 8542 21644
rect 3878 21564 3884 21616
rect 3936 21604 3942 21616
rect 4706 21604 4712 21616
rect 3936 21576 4712 21604
rect 3936 21564 3942 21576
rect 4706 21564 4712 21576
rect 4764 21604 4770 21616
rect 5718 21604 5724 21616
rect 4764 21576 5724 21604
rect 4764 21564 4770 21576
rect 5718 21564 5724 21576
rect 5776 21564 5782 21616
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 9125 21607 9183 21613
rect 9125 21604 9137 21607
rect 8996 21576 9137 21604
rect 8996 21564 9002 21576
rect 9125 21573 9137 21576
rect 9171 21573 9183 21607
rect 9674 21604 9680 21616
rect 9125 21567 9183 21573
rect 9140 21536 9168 21567
rect 9646 21564 9680 21604
rect 9732 21564 9738 21616
rect 10612 21604 10640 21644
rect 10686 21632 10692 21684
rect 10744 21672 10750 21684
rect 11057 21675 11115 21681
rect 11057 21672 11069 21675
rect 10744 21644 11069 21672
rect 10744 21632 10750 21644
rect 11057 21641 11069 21644
rect 11103 21641 11115 21675
rect 11057 21635 11115 21641
rect 12342 21632 12348 21684
rect 12400 21672 12406 21684
rect 12400 21644 16988 21672
rect 12400 21632 12406 21644
rect 14074 21607 14132 21613
rect 10612 21576 10732 21604
rect 9646 21536 9674 21564
rect 5552 21508 6960 21536
rect 9140 21508 9674 21536
rect 10704 21536 10732 21576
rect 14074 21573 14086 21607
rect 14120 21604 14132 21607
rect 14826 21604 14832 21616
rect 14120 21576 14832 21604
rect 14120 21573 14132 21576
rect 14074 21567 14132 21573
rect 14826 21564 14832 21576
rect 14884 21564 14890 21616
rect 16114 21564 16120 21616
rect 16172 21604 16178 21616
rect 16390 21604 16396 21616
rect 16172 21576 16396 21604
rect 16172 21564 16178 21576
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 12894 21536 12900 21548
rect 10704 21508 12900 21536
rect 1670 21468 1676 21480
rect 1631 21440 1676 21468
rect 1670 21428 1676 21440
rect 1728 21428 1734 21480
rect 2130 21468 2136 21480
rect 2091 21440 2136 21468
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3602 21468 3608 21480
rect 2823 21440 3608 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 4709 21471 4767 21477
rect 4709 21468 4721 21471
rect 4172 21440 4721 21468
rect 3044 21403 3102 21409
rect 3044 21369 3056 21403
rect 3090 21400 3102 21403
rect 3326 21400 3332 21412
rect 3090 21372 3332 21400
rect 3090 21369 3102 21372
rect 3044 21363 3102 21369
rect 3326 21360 3332 21372
rect 3384 21360 3390 21412
rect 4172 21344 4200 21440
rect 4709 21437 4721 21440
rect 4755 21437 4767 21471
rect 4709 21431 4767 21437
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5442 21468 5448 21480
rect 5399 21440 5448 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5442 21428 5448 21440
rect 5500 21428 5506 21480
rect 5552 21477 5580 21508
rect 6932 21480 6960 21508
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 14277 21539 14335 21545
rect 14277 21536 14289 21539
rect 13688 21508 14289 21536
rect 13688 21496 13694 21508
rect 14277 21505 14289 21508
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 15010 21496 15016 21548
rect 15068 21536 15074 21548
rect 15197 21539 15255 21545
rect 15197 21536 15209 21539
rect 15068 21508 15209 21536
rect 15068 21496 15074 21508
rect 15197 21505 15209 21508
rect 15243 21505 15255 21539
rect 16960 21536 16988 21644
rect 18230 21632 18236 21684
rect 18288 21672 18294 21684
rect 18325 21675 18383 21681
rect 18325 21672 18337 21675
rect 18288 21644 18337 21672
rect 18288 21632 18294 21644
rect 18325 21641 18337 21644
rect 18371 21672 18383 21675
rect 18414 21672 18420 21684
rect 18371 21644 18420 21672
rect 18371 21641 18383 21644
rect 18325 21635 18383 21641
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19242 21632 19248 21684
rect 19300 21672 19306 21684
rect 23014 21672 23020 21684
rect 19300 21644 22876 21672
rect 22975 21644 23020 21672
rect 19300 21632 19306 21644
rect 17034 21564 17040 21616
rect 17092 21604 17098 21616
rect 17494 21604 17500 21616
rect 17092 21576 17500 21604
rect 17092 21564 17098 21576
rect 17494 21564 17500 21576
rect 17552 21564 17558 21616
rect 17586 21564 17592 21616
rect 17644 21604 17650 21616
rect 17644 21576 18920 21604
rect 17644 21564 17650 21576
rect 16960 21508 18184 21536
rect 15197 21499 15255 21505
rect 5537 21471 5595 21477
rect 5537 21437 5549 21471
rect 5583 21437 5595 21471
rect 5718 21468 5724 21480
rect 5679 21440 5724 21468
rect 5537 21431 5595 21437
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 6362 21468 6368 21480
rect 5868 21440 6368 21468
rect 5868 21428 5874 21440
rect 6362 21428 6368 21440
rect 6420 21428 6426 21480
rect 6638 21428 6644 21480
rect 6696 21468 6702 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6696 21440 6837 21468
rect 6696 21428 6702 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 6914 21428 6920 21480
rect 6972 21428 6978 21480
rect 7092 21471 7150 21477
rect 7092 21437 7104 21471
rect 7138 21468 7150 21471
rect 7374 21468 7380 21480
rect 7138 21440 7380 21468
rect 7138 21437 7150 21440
rect 7092 21431 7150 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 8846 21468 8852 21480
rect 8807 21440 8852 21468
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 8941 21471 8999 21477
rect 8941 21437 8953 21471
rect 8987 21437 8999 21471
rect 9214 21468 9220 21480
rect 9175 21440 9220 21468
rect 8941 21431 8999 21437
rect 5629 21403 5687 21409
rect 5629 21369 5641 21403
rect 5675 21400 5687 21403
rect 7558 21400 7564 21412
rect 5675 21372 7564 21400
rect 5675 21369 5687 21372
rect 5629 21363 5687 21369
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 8294 21360 8300 21412
rect 8352 21400 8358 21412
rect 8956 21400 8984 21431
rect 9214 21428 9220 21440
rect 9272 21428 9278 21480
rect 9674 21468 9680 21480
rect 9635 21440 9680 21468
rect 9674 21428 9680 21440
rect 9732 21428 9738 21480
rect 9950 21477 9956 21480
rect 9944 21468 9956 21477
rect 9911 21440 9956 21468
rect 9944 21431 9956 21440
rect 9950 21428 9956 21431
rect 10008 21428 10014 21480
rect 12342 21468 12348 21480
rect 10051 21440 12348 21468
rect 10051 21400 10079 21440
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 12710 21468 12716 21480
rect 12575 21440 12716 21468
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 13265 21471 13323 21477
rect 13265 21437 13277 21471
rect 13311 21468 13323 21471
rect 13722 21468 13728 21480
rect 13311 21440 13728 21468
rect 13311 21437 13323 21440
rect 13265 21431 13323 21437
rect 13722 21428 13728 21440
rect 13780 21428 13786 21480
rect 14182 21477 14188 21480
rect 14139 21471 14188 21477
rect 14139 21437 14151 21471
rect 14185 21437 14188 21471
rect 14139 21431 14188 21437
rect 14182 21428 14188 21431
rect 14240 21428 14246 21480
rect 15105 21471 15163 21477
rect 15105 21437 15117 21471
rect 15151 21437 15163 21471
rect 15105 21431 15163 21437
rect 8352 21372 10079 21400
rect 13909 21403 13967 21409
rect 8352 21360 8358 21372
rect 13909 21369 13921 21403
rect 13955 21369 13967 21403
rect 15120 21400 15148 21431
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 15381 21471 15439 21477
rect 15381 21468 15393 21471
rect 15344 21440 15393 21468
rect 15344 21428 15350 21440
rect 15381 21437 15393 21440
rect 15427 21437 15439 21471
rect 15381 21431 15439 21437
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15841 21471 15899 21477
rect 15841 21468 15853 21471
rect 15528 21440 15853 21468
rect 15528 21428 15534 21440
rect 15841 21437 15853 21440
rect 15887 21468 15899 21471
rect 17034 21468 17040 21480
rect 15887 21440 17040 21468
rect 15887 21437 15899 21440
rect 15841 21431 15899 21437
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 18156 21477 18184 21508
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 18141 21471 18199 21477
rect 18141 21437 18153 21471
rect 18187 21468 18199 21471
rect 18230 21468 18236 21480
rect 18187 21440 18236 21468
rect 18187 21437 18199 21440
rect 18141 21431 18199 21437
rect 15930 21400 15936 21412
rect 15120 21372 15936 21400
rect 13909 21363 13967 21369
rect 1489 21335 1547 21341
rect 1489 21301 1501 21335
rect 1535 21332 1547 21335
rect 3786 21332 3792 21344
rect 1535 21304 3792 21332
rect 1535 21301 1547 21304
rect 1489 21295 1547 21301
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 4154 21332 4160 21344
rect 4115 21304 4160 21332
rect 4154 21292 4160 21304
rect 4212 21292 4218 21344
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 4890 21332 4896 21344
rect 4847 21304 4896 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 4890 21292 4896 21304
rect 4948 21292 4954 21344
rect 5902 21292 5908 21344
rect 5960 21332 5966 21344
rect 8665 21335 8723 21341
rect 5960 21304 6005 21332
rect 5960 21292 5966 21304
rect 8665 21301 8677 21335
rect 8711 21332 8723 21335
rect 9306 21332 9312 21344
rect 8711 21304 9312 21332
rect 8711 21301 8723 21304
rect 8665 21295 8723 21301
rect 9306 21292 9312 21304
rect 9364 21292 9370 21344
rect 9398 21292 9404 21344
rect 9456 21332 9462 21344
rect 10778 21332 10784 21344
rect 9456 21304 10784 21332
rect 9456 21292 9462 21304
rect 10778 21292 10784 21304
rect 10836 21332 10842 21344
rect 12618 21332 12624 21344
rect 10836 21304 12624 21332
rect 10836 21292 10842 21304
rect 12618 21292 12624 21304
rect 12676 21292 12682 21344
rect 12713 21335 12771 21341
rect 12713 21301 12725 21335
rect 12759 21332 12771 21335
rect 13262 21332 13268 21344
rect 12759 21304 13268 21332
rect 12759 21301 12771 21304
rect 12713 21295 12771 21301
rect 13262 21292 13268 21304
rect 13320 21292 13326 21344
rect 13357 21335 13415 21341
rect 13357 21301 13369 21335
rect 13403 21332 13415 21335
rect 13722 21332 13728 21344
rect 13403 21304 13728 21332
rect 13403 21301 13415 21304
rect 13357 21295 13415 21301
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 13924 21332 13952 21363
rect 15930 21360 15936 21372
rect 15988 21360 15994 21412
rect 18064 21400 18092 21431
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18417 21471 18475 21477
rect 18417 21437 18429 21471
rect 18463 21468 18475 21471
rect 18598 21468 18604 21480
rect 18463 21440 18604 21468
rect 18463 21437 18475 21440
rect 18417 21431 18475 21437
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 18892 21477 18920 21576
rect 18966 21564 18972 21616
rect 19024 21604 19030 21616
rect 19024 21576 19334 21604
rect 19024 21564 19030 21576
rect 19306 21536 19334 21576
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19306 21508 19533 21536
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 20956 21508 22094 21536
rect 20956 21496 20962 21508
rect 18877 21471 18935 21477
rect 18877 21437 18889 21471
rect 18923 21437 18935 21471
rect 18877 21431 18935 21437
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 19150 21468 19156 21480
rect 19024 21440 19156 21468
rect 19024 21428 19030 21440
rect 19150 21428 19156 21440
rect 19208 21428 19214 21480
rect 19788 21471 19846 21477
rect 19788 21437 19800 21471
rect 19834 21468 19846 21471
rect 20530 21468 20536 21480
rect 19834 21440 20536 21468
rect 19834 21437 19846 21440
rect 19788 21431 19846 21437
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 20622 21428 20628 21480
rect 20680 21468 20686 21480
rect 21361 21471 21419 21477
rect 21361 21468 21373 21471
rect 20680 21440 21373 21468
rect 20680 21428 20686 21440
rect 21361 21437 21373 21440
rect 21407 21437 21419 21471
rect 21361 21431 21419 21437
rect 21453 21403 21511 21409
rect 21453 21400 21465 21403
rect 18064 21372 21465 21400
rect 21453 21369 21465 21372
rect 21499 21369 21511 21403
rect 22066 21400 22094 21508
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 22848 21477 22876 21644
rect 23014 21632 23020 21644
rect 23072 21632 23078 21684
rect 24210 21672 24216 21684
rect 24171 21644 24216 21672
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 25406 21672 25412 21684
rect 25367 21644 25412 21672
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 23198 21564 23204 21616
rect 23256 21604 23262 21616
rect 23658 21604 23664 21616
rect 23256 21576 23664 21604
rect 23256 21564 23262 21576
rect 23658 21564 23664 21576
rect 23716 21604 23722 21616
rect 23934 21604 23940 21616
rect 23716 21576 23940 21604
rect 23716 21564 23722 21576
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 25682 21564 25688 21616
rect 25740 21604 25746 21616
rect 25740 21576 26372 21604
rect 25740 21564 25746 21576
rect 24578 21536 24584 21548
rect 23124 21508 24584 21536
rect 23124 21477 23152 21508
rect 24578 21496 24584 21508
rect 24636 21496 24642 21548
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22704 21440 22753 21468
rect 22704 21428 22710 21440
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 22833 21471 22891 21477
rect 22833 21437 22845 21471
rect 22879 21437 22891 21471
rect 22833 21431 22891 21437
rect 23109 21471 23167 21477
rect 23109 21437 23121 21471
rect 23155 21437 23167 21471
rect 23109 21431 23167 21437
rect 23566 21428 23572 21480
rect 23624 21468 23630 21480
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 23624 21440 23673 21468
rect 23624 21428 23630 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23934 21468 23940 21480
rect 23895 21440 23940 21468
rect 23661 21431 23719 21437
rect 23934 21428 23940 21440
rect 23992 21428 23998 21480
rect 24029 21471 24087 21477
rect 24029 21437 24041 21471
rect 24075 21468 24087 21471
rect 24302 21468 24308 21480
rect 24075 21440 24308 21468
rect 24075 21437 24087 21440
rect 24029 21431 24087 21437
rect 24302 21428 24308 21440
rect 24360 21428 24366 21480
rect 24486 21428 24492 21480
rect 24544 21468 24550 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 24544 21440 24685 21468
rect 24544 21428 24550 21440
rect 24673 21437 24685 21440
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 25317 21471 25375 21477
rect 25317 21437 25329 21471
rect 25363 21468 25375 21471
rect 25590 21468 25596 21480
rect 25363 21440 25596 21468
rect 25363 21437 25375 21440
rect 25317 21431 25375 21437
rect 25590 21428 25596 21440
rect 25648 21428 25654 21480
rect 26344 21477 26372 21576
rect 25961 21471 26019 21477
rect 25961 21437 25973 21471
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21437 26295 21471
rect 26237 21431 26295 21437
rect 26329 21471 26387 21477
rect 26329 21437 26341 21471
rect 26375 21437 26387 21471
rect 26329 21431 26387 21437
rect 23845 21403 23903 21409
rect 22066 21372 23796 21400
rect 21453 21363 21511 21369
rect 14274 21332 14280 21344
rect 13924 21304 14280 21332
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14553 21335 14611 21341
rect 14553 21301 14565 21335
rect 14599 21332 14611 21335
rect 15102 21332 15108 21344
rect 14599 21304 15108 21332
rect 14599 21301 14611 21304
rect 14553 21295 14611 21301
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 15194 21292 15200 21344
rect 15252 21332 15258 21344
rect 16114 21332 16120 21344
rect 15252 21304 16120 21332
rect 15252 21292 15258 21304
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 17865 21335 17923 21341
rect 17865 21301 17877 21335
rect 17911 21332 17923 21335
rect 18046 21332 18052 21344
rect 17911 21304 18052 21332
rect 17911 21301 17923 21304
rect 17865 21295 17923 21301
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 18598 21292 18604 21344
rect 18656 21332 18662 21344
rect 18969 21335 19027 21341
rect 18969 21332 18981 21335
rect 18656 21304 18981 21332
rect 18656 21292 18662 21304
rect 18969 21301 18981 21304
rect 19015 21301 19027 21335
rect 18969 21295 19027 21301
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 20254 21332 20260 21344
rect 19576 21304 20260 21332
rect 19576 21292 19582 21304
rect 20254 21292 20260 21304
rect 20312 21332 20318 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20312 21304 20913 21332
rect 20312 21292 20318 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 20901 21295 20959 21301
rect 22557 21335 22615 21341
rect 22557 21301 22569 21335
rect 22603 21332 22615 21335
rect 23106 21332 23112 21344
rect 22603 21304 23112 21332
rect 22603 21301 22615 21304
rect 22557 21295 22615 21301
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 23768 21332 23796 21372
rect 23845 21369 23857 21403
rect 23891 21400 23903 21403
rect 24210 21400 24216 21412
rect 23891 21372 24216 21400
rect 23891 21369 23903 21372
rect 23845 21363 23903 21369
rect 24210 21360 24216 21372
rect 24268 21400 24274 21412
rect 24762 21400 24768 21412
rect 24268 21372 24768 21400
rect 24268 21360 24274 21372
rect 24762 21360 24768 21372
rect 24820 21360 24826 21412
rect 25222 21360 25228 21412
rect 25280 21400 25286 21412
rect 25976 21400 26004 21431
rect 25280 21372 26004 21400
rect 26145 21403 26203 21409
rect 25280 21360 25286 21372
rect 26145 21369 26157 21403
rect 26191 21369 26203 21403
rect 26252 21400 26280 21431
rect 26970 21400 26976 21412
rect 26252 21372 26976 21400
rect 26145 21363 26203 21369
rect 25682 21332 25688 21344
rect 23768 21304 25688 21332
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 25774 21292 25780 21344
rect 25832 21332 25838 21344
rect 26160 21332 26188 21363
rect 26970 21360 26976 21372
rect 27028 21360 27034 21412
rect 26510 21332 26516 21344
rect 25832 21304 26188 21332
rect 26471 21304 26516 21332
rect 25832 21292 25838 21304
rect 26510 21292 26516 21304
rect 26568 21292 26574 21344
rect 1104 21242 28428 21264
rect 1104 21190 10090 21242
rect 10142 21190 10154 21242
rect 10206 21190 10218 21242
rect 10270 21190 10282 21242
rect 10334 21190 19198 21242
rect 19250 21190 19262 21242
rect 19314 21190 19326 21242
rect 19378 21190 19390 21242
rect 19442 21190 28428 21242
rect 1104 21168 28428 21190
rect 1946 21128 1952 21140
rect 1907 21100 1952 21128
rect 1946 21088 1952 21100
rect 2004 21088 2010 21140
rect 3326 21128 3332 21140
rect 3287 21100 3332 21128
rect 3326 21088 3332 21100
rect 3384 21088 3390 21140
rect 5994 21128 6000 21140
rect 4724 21100 6000 21128
rect 3053 21063 3111 21069
rect 3053 21029 3065 21063
rect 3099 21060 3111 21063
rect 4154 21060 4160 21072
rect 3099 21032 4160 21060
rect 3099 21029 3111 21032
rect 3053 21023 3111 21029
rect 4154 21020 4160 21032
rect 4212 21020 4218 21072
rect 1854 20992 1860 21004
rect 1815 20964 1860 20992
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20961 2835 20995
rect 2777 20955 2835 20961
rect 2961 20995 3019 21001
rect 2961 20961 2973 20995
rect 3007 20961 3019 20995
rect 2961 20955 3019 20961
rect 3145 20995 3203 21001
rect 3145 20961 3157 20995
rect 3191 20992 3203 20995
rect 3878 20992 3884 21004
rect 3191 20964 3884 20992
rect 3191 20961 3203 20964
rect 3145 20955 3203 20961
rect 2792 20788 2820 20955
rect 2976 20924 3004 20955
rect 3878 20952 3884 20964
rect 3936 20952 3942 21004
rect 4724 21001 4752 21100
rect 5994 21088 6000 21100
rect 6052 21088 6058 21140
rect 6362 21088 6368 21140
rect 6420 21128 6426 21140
rect 9398 21128 9404 21140
rect 6420 21100 9404 21128
rect 6420 21088 6426 21100
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 9674 21088 9680 21140
rect 9732 21128 9738 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 9732 21100 10333 21128
rect 9732 21088 9738 21100
rect 10321 21097 10333 21100
rect 10367 21128 10379 21131
rect 10778 21128 10784 21140
rect 10367 21100 10784 21128
rect 10367 21097 10379 21100
rect 10321 21091 10379 21097
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 10870 21088 10876 21140
rect 10928 21128 10934 21140
rect 11793 21131 11851 21137
rect 11793 21128 11805 21131
rect 10928 21100 11805 21128
rect 10928 21088 10934 21100
rect 11793 21097 11805 21100
rect 11839 21128 11851 21131
rect 11839 21100 19334 21128
rect 11839 21097 11851 21100
rect 11793 21091 11851 21097
rect 5810 21060 5816 21072
rect 5000 21032 5816 21060
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20961 4767 20995
rect 4890 20992 4896 21004
rect 4851 20964 4896 20992
rect 4709 20955 4767 20961
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 5000 21001 5028 21032
rect 5810 21020 5816 21032
rect 5868 21020 5874 21072
rect 5902 21020 5908 21072
rect 5960 21060 5966 21072
rect 6150 21063 6208 21069
rect 6150 21060 6162 21063
rect 5960 21032 6162 21060
rect 5960 21020 5966 21032
rect 6150 21029 6162 21032
rect 6196 21029 6208 21063
rect 6150 21023 6208 21029
rect 6730 21020 6736 21072
rect 6788 21060 6794 21072
rect 6788 21032 9628 21060
rect 6788 21020 6794 21032
rect 4985 20995 5043 21001
rect 4985 20961 4997 20995
rect 5031 20961 5043 20995
rect 5258 20992 5264 21004
rect 5219 20964 5264 20992
rect 4985 20955 5043 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5445 20995 5503 21001
rect 5445 20961 5457 20995
rect 5491 20992 5503 20995
rect 7926 20992 7932 21004
rect 5491 20964 7932 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 8205 20995 8263 21001
rect 8205 20961 8217 20995
rect 8251 20961 8263 20995
rect 8205 20955 8263 20961
rect 3050 20924 3056 20936
rect 2976 20896 3056 20924
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 5077 20927 5135 20933
rect 5077 20893 5089 20927
rect 5123 20924 5135 20927
rect 5810 20924 5816 20936
rect 5123 20896 5816 20924
rect 5123 20893 5135 20896
rect 5077 20887 5135 20893
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 4246 20788 4252 20800
rect 2792 20760 4252 20788
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 5920 20788 5948 20887
rect 8220 20856 8248 20955
rect 8294 20952 8300 21004
rect 8352 20992 8358 21004
rect 8573 20995 8631 21001
rect 8352 20964 8397 20992
rect 8352 20952 8358 20964
rect 8573 20961 8585 20995
rect 8619 20992 8631 20995
rect 8662 20992 8668 21004
rect 8619 20964 8668 20992
rect 8619 20961 8631 20964
rect 8573 20955 8631 20961
rect 8662 20952 8668 20964
rect 8720 20952 8726 21004
rect 9490 20992 9496 21004
rect 9451 20964 9496 20992
rect 9490 20952 9496 20964
rect 9548 20952 9554 21004
rect 9600 20992 9628 21032
rect 10410 21020 10416 21072
rect 10468 21060 10474 21072
rect 10658 21063 10716 21069
rect 10658 21060 10670 21063
rect 10468 21032 10670 21060
rect 10468 21020 10474 21032
rect 10658 21029 10670 21032
rect 10704 21029 10716 21063
rect 10658 21023 10716 21029
rect 12437 21063 12495 21069
rect 12437 21029 12449 21063
rect 12483 21060 12495 21063
rect 13817 21063 13875 21069
rect 12483 21032 13768 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 12618 20992 12624 21004
rect 9600 20964 12434 20992
rect 12579 20964 12624 20992
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20924 10379 20927
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 10367 20896 10425 20924
rect 10367 20893 10379 20896
rect 10321 20887 10379 20893
rect 10413 20893 10425 20896
rect 10459 20893 10471 20927
rect 12406 20924 12434 20964
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 13081 20995 13139 21001
rect 13081 20961 13093 20995
rect 13127 20992 13139 20995
rect 13354 20992 13360 21004
rect 13127 20964 13360 20992
rect 13127 20961 13139 20964
rect 13081 20955 13139 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 13740 20992 13768 21032
rect 13817 21029 13829 21063
rect 13863 21060 13875 21063
rect 15930 21060 15936 21072
rect 13863 21032 15936 21060
rect 13863 21029 13875 21032
rect 13817 21023 13875 21029
rect 15930 21020 15936 21032
rect 15988 21020 15994 21072
rect 16025 21063 16083 21069
rect 16025 21029 16037 21063
rect 16071 21060 16083 21063
rect 17126 21060 17132 21072
rect 16071 21032 17132 21060
rect 16071 21029 16083 21032
rect 16025 21023 16083 21029
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 17405 21063 17463 21069
rect 17405 21029 17417 21063
rect 17451 21060 17463 21063
rect 17678 21060 17684 21072
rect 17451 21032 17684 21060
rect 17451 21029 17463 21032
rect 17405 21023 17463 21029
rect 17678 21020 17684 21032
rect 17736 21020 17742 21072
rect 19306 21060 19334 21100
rect 20070 21088 20076 21140
rect 20128 21128 20134 21140
rect 20165 21131 20223 21137
rect 20165 21128 20177 21131
rect 20128 21100 20177 21128
rect 20128 21088 20134 21100
rect 20165 21097 20177 21100
rect 20211 21097 20223 21131
rect 20165 21091 20223 21097
rect 21913 21131 21971 21137
rect 21913 21097 21925 21131
rect 21959 21128 21971 21131
rect 22462 21128 22468 21140
rect 21959 21100 22468 21128
rect 21959 21097 21971 21100
rect 21913 21091 21971 21097
rect 22462 21088 22468 21100
rect 22520 21088 22526 21140
rect 22646 21128 22652 21140
rect 22607 21100 22652 21128
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 24394 21128 24400 21140
rect 23216 21100 24400 21128
rect 20990 21060 20996 21072
rect 19306 21032 20996 21060
rect 20990 21020 20996 21032
rect 21048 21020 21054 21072
rect 21729 21063 21787 21069
rect 21729 21029 21741 21063
rect 21775 21060 21787 21063
rect 23014 21060 23020 21072
rect 21775 21032 23020 21060
rect 21775 21029 21787 21032
rect 21729 21023 21787 21029
rect 23014 21020 23020 21032
rect 23072 21020 23078 21072
rect 14458 20992 14464 21004
rect 13740 20964 14464 20992
rect 14458 20952 14464 20964
rect 14516 20992 14522 21004
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 14516 20964 14749 20992
rect 14516 20952 14522 20964
rect 14737 20961 14749 20964
rect 14783 20961 14795 20995
rect 14737 20955 14795 20961
rect 14826 20952 14832 21004
rect 14884 21001 14890 21004
rect 14884 20995 14942 21001
rect 14884 20961 14896 20995
rect 14930 20961 14942 20995
rect 14884 20955 14942 20961
rect 14884 20952 14890 20955
rect 15194 20952 15200 21004
rect 15252 20992 15258 21004
rect 15470 20992 15476 21004
rect 15252 20964 15476 20992
rect 15252 20952 15258 20964
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 17034 20952 17040 21004
rect 17092 20992 17098 21004
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 17092 20964 17233 20992
rect 17092 20952 17098 20964
rect 17221 20961 17233 20964
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20961 18199 20995
rect 18141 20955 18199 20961
rect 13449 20927 13507 20933
rect 12406 20896 13216 20924
rect 10413 20887 10471 20893
rect 8294 20856 8300 20868
rect 8220 20828 8300 20856
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 13188 20856 13216 20896
rect 13449 20893 13461 20927
rect 13495 20924 13507 20927
rect 13630 20924 13636 20936
rect 13495 20896 13636 20924
rect 13495 20893 13507 20896
rect 13449 20887 13507 20893
rect 13630 20884 13636 20896
rect 13688 20884 13694 20936
rect 13722 20884 13728 20936
rect 13780 20924 13786 20936
rect 15102 20924 15108 20936
rect 13780 20896 14964 20924
rect 15063 20896 15108 20924
rect 13780 20884 13786 20896
rect 13246 20859 13304 20865
rect 13246 20856 13258 20859
rect 13188 20828 13258 20856
rect 13246 20825 13258 20828
rect 13292 20856 13304 20859
rect 14826 20856 14832 20868
rect 13292 20828 14832 20856
rect 13292 20825 13304 20828
rect 13246 20819 13304 20825
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 14936 20856 14964 20896
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 17310 20924 17316 20936
rect 15212 20896 17316 20924
rect 15212 20856 15240 20896
rect 17310 20884 17316 20896
rect 17368 20884 17374 20936
rect 18156 20924 18184 20955
rect 18230 20952 18236 21004
rect 18288 20992 18294 21004
rect 18506 20992 18512 21004
rect 18288 20964 18333 20992
rect 18467 20964 18512 20992
rect 18288 20952 18294 20964
rect 18506 20952 18512 20964
rect 18564 20952 18570 21004
rect 18690 20952 18696 21004
rect 18748 20992 18754 21004
rect 18748 20964 19748 20992
rect 18748 20952 18754 20964
rect 19610 20924 19616 20936
rect 18156 20896 19616 20924
rect 19610 20884 19616 20896
rect 19668 20884 19674 20936
rect 19720 20924 19748 20964
rect 19978 20952 19984 21004
rect 20036 20992 20042 21004
rect 20073 20995 20131 21001
rect 20073 20992 20085 20995
rect 20036 20964 20085 20992
rect 20036 20952 20042 20964
rect 20073 20961 20085 20964
rect 20119 20992 20131 20995
rect 20438 20992 20444 21004
rect 20119 20964 20444 20992
rect 20119 20961 20131 20964
rect 20073 20955 20131 20961
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 20714 20992 20720 21004
rect 20675 20964 20720 20992
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 21818 20992 21824 21004
rect 21779 20964 21824 20992
rect 21818 20952 21824 20964
rect 21876 20952 21882 21004
rect 22554 20992 22560 21004
rect 22515 20964 22560 20992
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23216 21001 23244 21100
rect 24394 21088 24400 21100
rect 24452 21088 24458 21140
rect 25869 21131 25927 21137
rect 25869 21097 25881 21131
rect 25915 21097 25927 21131
rect 25869 21091 25927 21097
rect 25501 21063 25559 21069
rect 25501 21060 25513 21063
rect 25424 21032 25513 21060
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20961 23259 20995
rect 23201 20955 23259 20961
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24578 20992 24584 21004
rect 23891 20964 24584 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24578 20952 24584 20964
rect 24636 20952 24642 21004
rect 25222 20952 25228 21004
rect 25280 20992 25286 21004
rect 25317 20995 25375 21001
rect 25317 20992 25329 20995
rect 25280 20964 25329 20992
rect 25280 20952 25286 20964
rect 25317 20961 25329 20964
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 25332 20924 25360 20955
rect 19720 20896 25360 20924
rect 14936 20828 15240 20856
rect 15562 20816 15568 20868
rect 15620 20856 15626 20868
rect 16209 20859 16267 20865
rect 16209 20856 16221 20859
rect 15620 20828 16221 20856
rect 15620 20816 15626 20828
rect 16209 20825 16221 20828
rect 16255 20856 16267 20859
rect 18414 20856 18420 20868
rect 16255 20828 18092 20856
rect 18375 20828 18420 20856
rect 16255 20825 16267 20828
rect 16209 20819 16267 20825
rect 6178 20788 6184 20800
rect 5920 20760 6184 20788
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 7285 20791 7343 20797
rect 7285 20757 7297 20791
rect 7331 20788 7343 20791
rect 7558 20788 7564 20800
rect 7331 20760 7564 20788
rect 7331 20757 7343 20760
rect 7285 20751 7343 20757
rect 7558 20748 7564 20760
rect 7616 20748 7622 20800
rect 8021 20791 8079 20797
rect 8021 20757 8033 20791
rect 8067 20788 8079 20791
rect 8386 20788 8392 20800
rect 8067 20760 8392 20788
rect 8067 20757 8079 20760
rect 8021 20751 8079 20757
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 8481 20791 8539 20797
rect 8481 20757 8493 20791
rect 8527 20788 8539 20791
rect 8938 20788 8944 20800
rect 8527 20760 8944 20788
rect 8527 20757 8539 20760
rect 8481 20751 8539 20757
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20788 9643 20791
rect 10686 20788 10692 20800
rect 9631 20760 10692 20788
rect 9631 20757 9643 20760
rect 9585 20751 9643 20757
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 12250 20748 12256 20800
rect 12308 20788 12314 20800
rect 13357 20791 13415 20797
rect 13357 20788 13369 20791
rect 12308 20760 13369 20788
rect 12308 20748 12314 20760
rect 13357 20757 13369 20760
rect 13403 20788 13415 20791
rect 14182 20788 14188 20800
rect 13403 20760 14188 20788
rect 13403 20757 13415 20760
rect 13357 20751 13415 20757
rect 14182 20748 14188 20760
rect 14240 20788 14246 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14240 20760 15025 20788
rect 14240 20748 14246 20760
rect 15013 20757 15025 20760
rect 15059 20757 15071 20791
rect 15378 20788 15384 20800
rect 15339 20760 15384 20788
rect 15013 20751 15071 20757
rect 15378 20748 15384 20760
rect 15436 20788 15442 20800
rect 15838 20788 15844 20800
rect 15436 20760 15844 20788
rect 15436 20748 15442 20760
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 17770 20748 17776 20800
rect 17828 20788 17834 20800
rect 17957 20791 18015 20797
rect 17957 20788 17969 20791
rect 17828 20760 17969 20788
rect 17828 20748 17834 20760
rect 17957 20757 17969 20760
rect 18003 20757 18015 20791
rect 18064 20788 18092 20828
rect 18414 20816 18420 20828
rect 18472 20816 18478 20868
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 20809 20859 20867 20865
rect 20809 20856 20821 20859
rect 19392 20828 20821 20856
rect 19392 20816 19398 20828
rect 20809 20825 20821 20828
rect 20855 20825 20867 20859
rect 20809 20819 20867 20825
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 22462 20856 22468 20868
rect 21324 20828 22468 20856
rect 21324 20816 21330 20828
rect 22462 20816 22468 20828
rect 22520 20856 22526 20868
rect 25424 20856 25452 21032
rect 25501 21029 25513 21032
rect 25547 21029 25559 21063
rect 25884 21060 25912 21091
rect 26574 21063 26632 21069
rect 26574 21060 26586 21063
rect 25884 21032 26586 21060
rect 25501 21023 25559 21029
rect 26574 21029 26586 21032
rect 26620 21029 26632 21063
rect 26574 21023 26632 21029
rect 25590 20992 25596 21004
rect 25503 20964 25596 20992
rect 25590 20952 25596 20964
rect 25648 20952 25654 21004
rect 25682 20952 25688 21004
rect 25740 20992 25746 21004
rect 25740 20964 25785 20992
rect 25740 20952 25746 20964
rect 26050 20952 26056 21004
rect 26108 20992 26114 21004
rect 26329 20995 26387 21001
rect 26329 20992 26341 20995
rect 26108 20964 26341 20992
rect 26108 20952 26114 20964
rect 26329 20961 26341 20964
rect 26375 20961 26387 20995
rect 26329 20955 26387 20961
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 27338 20992 27344 21004
rect 27120 20964 27344 20992
rect 27120 20952 27126 20964
rect 27338 20952 27344 20964
rect 27396 20952 27402 21004
rect 22520 20828 25452 20856
rect 22520 20816 22526 20828
rect 21729 20791 21787 20797
rect 21729 20788 21741 20791
rect 18064 20760 21741 20788
rect 17957 20751 18015 20757
rect 21729 20757 21741 20760
rect 21775 20757 21787 20791
rect 21729 20751 21787 20757
rect 23293 20791 23351 20797
rect 23293 20757 23305 20791
rect 23339 20788 23351 20791
rect 23474 20788 23480 20800
rect 23339 20760 23480 20788
rect 23339 20757 23351 20760
rect 23293 20751 23351 20757
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 23937 20791 23995 20797
rect 23937 20757 23949 20791
rect 23983 20788 23995 20791
rect 24118 20788 24124 20800
rect 23983 20760 24124 20788
rect 23983 20757 23995 20760
rect 23937 20751 23995 20757
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 25608 20788 25636 20952
rect 27338 20788 27344 20800
rect 25608 20760 27344 20788
rect 27338 20748 27344 20760
rect 27396 20788 27402 20800
rect 27709 20791 27767 20797
rect 27709 20788 27721 20791
rect 27396 20760 27721 20788
rect 27396 20748 27402 20760
rect 27709 20757 27721 20760
rect 27755 20757 27767 20791
rect 27709 20751 27767 20757
rect 1104 20698 28428 20720
rect 1104 20646 5536 20698
rect 5588 20646 5600 20698
rect 5652 20646 5664 20698
rect 5716 20646 5728 20698
rect 5780 20646 14644 20698
rect 14696 20646 14708 20698
rect 14760 20646 14772 20698
rect 14824 20646 14836 20698
rect 14888 20646 23752 20698
rect 23804 20646 23816 20698
rect 23868 20646 23880 20698
rect 23932 20646 23944 20698
rect 23996 20646 28428 20698
rect 1104 20624 28428 20646
rect 3605 20587 3663 20593
rect 3605 20553 3617 20587
rect 3651 20584 3663 20587
rect 5258 20584 5264 20596
rect 3651 20556 5264 20584
rect 3651 20553 3663 20556
rect 3605 20547 3663 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 5902 20544 5908 20596
rect 5960 20584 5966 20596
rect 7098 20584 7104 20596
rect 5960 20556 7104 20584
rect 5960 20544 5966 20556
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 8570 20584 8576 20596
rect 8483 20556 8576 20584
rect 8570 20544 8576 20556
rect 8628 20584 8634 20596
rect 9490 20584 9496 20596
rect 8628 20556 9496 20584
rect 8628 20544 8634 20556
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 12342 20544 12348 20596
rect 12400 20584 12406 20596
rect 12437 20587 12495 20593
rect 12437 20584 12449 20587
rect 12400 20556 12449 20584
rect 12400 20544 12406 20556
rect 12437 20553 12449 20556
rect 12483 20553 12495 20587
rect 12437 20547 12495 20553
rect 14182 20544 14188 20596
rect 14240 20584 14246 20596
rect 15102 20584 15108 20596
rect 14240 20556 15108 20584
rect 14240 20544 14246 20556
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 17497 20587 17555 20593
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 18414 20584 18420 20596
rect 17543 20556 18420 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 18414 20544 18420 20556
rect 18472 20544 18478 20596
rect 19610 20584 19616 20596
rect 19571 20556 19616 20584
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 25498 20584 25504 20596
rect 22066 20556 25504 20584
rect 10689 20519 10747 20525
rect 10689 20485 10701 20519
rect 10735 20516 10747 20519
rect 10962 20516 10968 20528
rect 10735 20488 10968 20516
rect 10735 20485 10747 20488
rect 10689 20479 10747 20485
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 13262 20476 13268 20528
rect 13320 20516 13326 20528
rect 13863 20519 13921 20525
rect 13863 20516 13875 20519
rect 13320 20488 13875 20516
rect 13320 20476 13326 20488
rect 13863 20485 13875 20488
rect 13909 20485 13921 20519
rect 13863 20479 13921 20485
rect 14001 20519 14059 20525
rect 14001 20485 14013 20519
rect 14047 20516 14059 20519
rect 16117 20519 16175 20525
rect 14047 20488 15047 20516
rect 14047 20485 14059 20488
rect 14001 20479 14059 20485
rect 6638 20408 6644 20460
rect 6696 20448 6702 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 6696 20420 7205 20448
rect 6696 20408 6702 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 10502 20448 10508 20460
rect 7193 20411 7251 20417
rect 10152 20420 10508 20448
rect 1578 20380 1584 20392
rect 1539 20352 1584 20380
rect 1578 20340 1584 20352
rect 1636 20340 1642 20392
rect 3513 20383 3571 20389
rect 3513 20349 3525 20383
rect 3559 20349 3571 20383
rect 3513 20343 3571 20349
rect 1848 20315 1906 20321
rect 1848 20281 1860 20315
rect 1894 20312 1906 20315
rect 2866 20312 2872 20324
rect 1894 20284 2872 20312
rect 1894 20281 1906 20284
rect 1848 20275 1906 20281
rect 2866 20272 2872 20284
rect 2924 20272 2930 20324
rect 2682 20204 2688 20256
rect 2740 20244 2746 20256
rect 2961 20247 3019 20253
rect 2961 20244 2973 20247
rect 2740 20216 2973 20244
rect 2740 20204 2746 20216
rect 2961 20213 2973 20216
rect 3007 20244 3019 20247
rect 3528 20244 3556 20343
rect 3602 20340 3608 20392
rect 3660 20380 3666 20392
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 3660 20352 4261 20380
rect 3660 20340 3666 20352
rect 4249 20349 4261 20352
rect 4295 20380 4307 20383
rect 6656 20380 6684 20408
rect 9306 20380 9312 20392
rect 4295 20352 6684 20380
rect 9267 20352 9312 20380
rect 4295 20349 4307 20352
rect 4249 20343 4307 20349
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 10152 20389 10180 20420
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10778 20448 10784 20460
rect 10739 20420 10784 20448
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 14090 20448 14096 20460
rect 14051 20420 14096 20448
rect 14090 20408 14096 20420
rect 14148 20448 14154 20460
rect 15019 20448 15047 20488
rect 16117 20485 16129 20519
rect 16163 20516 16175 20519
rect 22066 20516 22094 20556
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 16163 20488 22094 20516
rect 23845 20519 23903 20525
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 23845 20485 23857 20519
rect 23891 20516 23903 20519
rect 24762 20516 24768 20528
rect 23891 20488 24768 20516
rect 23891 20485 23903 20488
rect 23845 20479 23903 20485
rect 24762 20476 24768 20488
rect 24820 20476 24826 20528
rect 15746 20448 15752 20460
rect 14148 20420 14964 20448
rect 15019 20420 15752 20448
rect 14148 20408 14154 20420
rect 10137 20383 10195 20389
rect 10137 20349 10149 20383
rect 10183 20349 10195 20383
rect 10137 20343 10195 20349
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10410 20380 10416 20392
rect 10275 20352 10416 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10597 20383 10655 20389
rect 10597 20349 10609 20383
rect 10643 20349 10655 20383
rect 10597 20343 10655 20349
rect 4516 20315 4574 20321
rect 4516 20281 4528 20315
rect 4562 20312 4574 20315
rect 5810 20312 5816 20324
rect 4562 20284 5816 20312
rect 4562 20281 4574 20284
rect 4516 20275 4574 20281
rect 5810 20272 5816 20284
rect 5868 20272 5874 20324
rect 7466 20321 7472 20324
rect 7460 20275 7472 20321
rect 7524 20312 7530 20324
rect 7524 20284 7560 20312
rect 7466 20272 7472 20275
rect 7524 20272 7530 20284
rect 10502 20272 10508 20324
rect 10560 20312 10566 20324
rect 10612 20312 10640 20343
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 11238 20380 11244 20392
rect 11112 20352 11244 20380
rect 11112 20340 11118 20352
rect 11238 20340 11244 20352
rect 11296 20380 11302 20392
rect 13078 20380 13084 20392
rect 11296 20352 13084 20380
rect 11296 20340 11302 20352
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 13265 20383 13323 20389
rect 13265 20349 13277 20383
rect 13311 20380 13323 20383
rect 14936 20380 14964 20420
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 18966 20448 18972 20460
rect 18892 20420 18972 20448
rect 15102 20380 15108 20392
rect 13311 20352 13860 20380
rect 14936 20352 15108 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 10560 20284 10640 20312
rect 12345 20315 12403 20321
rect 10560 20272 10566 20284
rect 12345 20281 12357 20315
rect 12391 20281 12403 20315
rect 13722 20312 13728 20324
rect 13683 20284 13728 20312
rect 12345 20275 12403 20281
rect 3007 20216 3556 20244
rect 3007 20213 3019 20216
rect 2961 20207 3019 20213
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5629 20247 5687 20253
rect 5629 20244 5641 20247
rect 5592 20216 5641 20244
rect 5592 20204 5598 20216
rect 5629 20213 5641 20216
rect 5675 20213 5687 20247
rect 12360 20244 12388 20275
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 13832 20312 13860 20352
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 15286 20380 15292 20392
rect 15247 20352 15292 20380
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 15841 20383 15899 20389
rect 15841 20349 15853 20383
rect 15887 20380 15899 20383
rect 15930 20380 15936 20392
rect 15887 20352 15936 20380
rect 15887 20349 15899 20352
rect 15841 20343 15899 20349
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 18230 20340 18236 20392
rect 18288 20380 18294 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18288 20352 18521 20380
rect 18288 20340 18294 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 18690 20340 18696 20392
rect 18748 20380 18754 20392
rect 18892 20389 18920 20420
rect 18966 20408 18972 20420
rect 19024 20448 19030 20460
rect 23474 20448 23480 20460
rect 19024 20420 22094 20448
rect 23435 20420 23480 20448
rect 19024 20408 19030 20420
rect 18877 20383 18935 20389
rect 18877 20380 18889 20383
rect 18748 20352 18889 20380
rect 18748 20340 18754 20352
rect 18877 20349 18889 20352
rect 18923 20349 18935 20383
rect 18877 20343 18935 20349
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20380 19119 20383
rect 19334 20380 19340 20392
rect 19107 20352 19340 20380
rect 19107 20349 19119 20352
rect 19061 20343 19119 20349
rect 19334 20340 19340 20352
rect 19392 20340 19398 20392
rect 19518 20380 19524 20392
rect 19479 20352 19524 20380
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 20622 20380 20628 20392
rect 20583 20352 20628 20380
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20732 20352 21005 20380
rect 17218 20312 17224 20324
rect 13832 20284 17224 20312
rect 17218 20272 17224 20284
rect 17276 20312 17282 20324
rect 17405 20315 17463 20321
rect 17405 20312 17417 20315
rect 17276 20284 17417 20312
rect 17276 20272 17282 20284
rect 17405 20281 17417 20284
rect 17451 20281 17463 20315
rect 17405 20275 17463 20281
rect 18141 20315 18199 20321
rect 18141 20281 18153 20315
rect 18187 20312 18199 20315
rect 20070 20312 20076 20324
rect 18187 20284 20076 20312
rect 18187 20281 18199 20284
rect 18141 20275 18199 20281
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 20346 20272 20352 20324
rect 20404 20312 20410 20324
rect 20732 20312 20760 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 20993 20343 21051 20349
rect 20404 20284 20760 20312
rect 20809 20315 20867 20321
rect 20404 20272 20410 20284
rect 20809 20281 20821 20315
rect 20855 20281 20867 20315
rect 20809 20275 20867 20281
rect 20901 20315 20959 20321
rect 20901 20281 20913 20315
rect 20947 20312 20959 20315
rect 21818 20312 21824 20324
rect 20947 20284 21824 20312
rect 20947 20281 20959 20284
rect 20901 20275 20959 20281
rect 14274 20244 14280 20256
rect 12360 20216 14280 20244
rect 5629 20207 5687 20213
rect 14274 20204 14280 20216
rect 14332 20244 14338 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 14332 20216 14381 20244
rect 14332 20204 14338 20216
rect 14369 20213 14381 20216
rect 14415 20213 14427 20247
rect 14369 20207 14427 20213
rect 18782 20204 18788 20256
rect 18840 20244 18846 20256
rect 20824 20244 20852 20275
rect 21818 20272 21824 20284
rect 21876 20272 21882 20324
rect 22066 20312 22094 20420
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 23106 20380 23112 20392
rect 23067 20352 23112 20380
rect 23106 20340 23112 20352
rect 23164 20340 23170 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23569 20383 23627 20389
rect 23569 20380 23581 20383
rect 23348 20352 23581 20380
rect 23348 20340 23354 20352
rect 23569 20349 23581 20352
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 23937 20383 23995 20389
rect 23937 20349 23949 20383
rect 23983 20349 23995 20383
rect 24118 20380 24124 20392
rect 24079 20352 24124 20380
rect 23937 20343 23995 20349
rect 23382 20312 23388 20324
rect 22066 20284 23388 20312
rect 23382 20272 23388 20284
rect 23440 20312 23446 20324
rect 23952 20312 23980 20343
rect 24118 20340 24124 20352
rect 24176 20340 24182 20392
rect 24854 20380 24860 20392
rect 24815 20352 24860 20380
rect 24854 20340 24860 20352
rect 24912 20340 24918 20392
rect 25501 20383 25559 20389
rect 25501 20349 25513 20383
rect 25547 20349 25559 20383
rect 25501 20343 25559 20349
rect 25768 20383 25826 20389
rect 25768 20349 25780 20383
rect 25814 20380 25826 20383
rect 26510 20380 26516 20392
rect 25814 20352 26516 20380
rect 25814 20349 25826 20352
rect 25768 20343 25826 20349
rect 23440 20284 23980 20312
rect 25041 20315 25099 20321
rect 23440 20272 23446 20284
rect 25041 20281 25053 20315
rect 25087 20312 25099 20315
rect 25130 20312 25136 20324
rect 25087 20284 25136 20312
rect 25087 20281 25099 20284
rect 25041 20275 25099 20281
rect 25130 20272 25136 20284
rect 25188 20272 25194 20324
rect 25516 20312 25544 20343
rect 26510 20340 26516 20352
rect 26568 20340 26574 20392
rect 25516 20284 25820 20312
rect 25792 20256 25820 20284
rect 21174 20244 21180 20256
rect 18840 20216 20852 20244
rect 21135 20216 21180 20244
rect 18840 20204 18846 20216
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 25774 20204 25780 20256
rect 25832 20204 25838 20256
rect 26881 20247 26939 20253
rect 26881 20213 26893 20247
rect 26927 20244 26939 20247
rect 26970 20244 26976 20256
rect 26927 20216 26976 20244
rect 26927 20213 26939 20216
rect 26881 20207 26939 20213
rect 26970 20204 26976 20216
rect 27028 20204 27034 20256
rect 1104 20154 28428 20176
rect 1104 20102 10090 20154
rect 10142 20102 10154 20154
rect 10206 20102 10218 20154
rect 10270 20102 10282 20154
rect 10334 20102 19198 20154
rect 19250 20102 19262 20154
rect 19314 20102 19326 20154
rect 19378 20102 19390 20154
rect 19442 20102 28428 20154
rect 1104 20080 28428 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2924 20012 2973 20040
rect 2924 20000 2930 20012
rect 2961 20009 2973 20012
rect 3007 20009 3019 20043
rect 5810 20040 5816 20052
rect 5771 20012 5816 20040
rect 2961 20003 3019 20009
rect 5810 20000 5816 20012
rect 5868 20000 5874 20052
rect 6270 20040 6276 20052
rect 6231 20012 6276 20040
rect 6270 20000 6276 20012
rect 6328 20040 6334 20052
rect 6730 20040 6736 20052
rect 6328 20012 6736 20040
rect 6328 20000 6334 20012
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 7466 20040 7472 20052
rect 7427 20012 7472 20040
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 8294 20040 8300 20052
rect 8255 20012 8300 20040
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 10502 20040 10508 20052
rect 9732 20012 10508 20040
rect 9732 20000 9738 20012
rect 10502 20000 10508 20012
rect 10560 20040 10566 20052
rect 10560 20012 10824 20040
rect 10560 20000 10566 20012
rect 2593 19975 2651 19981
rect 2593 19941 2605 19975
rect 2639 19972 2651 19975
rect 3050 19972 3056 19984
rect 2639 19944 3056 19972
rect 2639 19941 2651 19944
rect 2593 19935 2651 19941
rect 3050 19932 3056 19944
rect 3108 19972 3114 19984
rect 5534 19972 5540 19984
rect 3108 19944 5396 19972
rect 5495 19944 5540 19972
rect 3108 19932 3114 19944
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 2222 19904 2228 19916
rect 1811 19876 2228 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 2406 19904 2412 19916
rect 2367 19876 2412 19904
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 2682 19904 2688 19916
rect 2595 19876 2688 19904
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3970 19904 3976 19916
rect 2823 19876 3976 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3970 19864 3976 19876
rect 4028 19864 4034 19916
rect 5261 19907 5319 19913
rect 5261 19873 5273 19907
rect 5307 19873 5319 19907
rect 5368 19904 5396 19944
rect 5534 19932 5540 19944
rect 5592 19972 5598 19984
rect 5902 19972 5908 19984
rect 5592 19944 5908 19972
rect 5592 19932 5598 19944
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 6546 19972 6552 19984
rect 6380 19944 6552 19972
rect 5442 19904 5448 19916
rect 5368 19876 5448 19904
rect 5261 19867 5319 19873
rect 1670 19796 1676 19848
rect 1728 19836 1734 19848
rect 2700 19836 2728 19864
rect 1728 19808 2728 19836
rect 5276 19836 5304 19867
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 5994 19904 6000 19916
rect 5675 19876 6000 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 5994 19864 6000 19876
rect 6052 19904 6058 19916
rect 6380 19904 6408 19944
rect 6546 19932 6552 19944
rect 6604 19932 6610 19984
rect 7006 19932 7012 19984
rect 7064 19972 7070 19984
rect 7101 19975 7159 19981
rect 7101 19972 7113 19975
rect 7064 19944 7113 19972
rect 7064 19932 7070 19944
rect 7101 19941 7113 19944
rect 7147 19941 7159 19975
rect 7101 19935 7159 19941
rect 7193 19975 7251 19981
rect 7193 19941 7205 19975
rect 7239 19972 7251 19975
rect 8570 19972 8576 19984
rect 7239 19944 8576 19972
rect 7239 19941 7251 19944
rect 7193 19935 7251 19941
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 6052 19876 6408 19904
rect 6457 19907 6515 19913
rect 6052 19864 6058 19876
rect 6457 19873 6469 19907
rect 6503 19873 6515 19907
rect 6914 19904 6920 19916
rect 6875 19876 6920 19904
rect 6457 19867 6515 19873
rect 6362 19836 6368 19848
rect 5276 19808 6368 19836
rect 1728 19796 1734 19808
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 6472 19836 6500 19867
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 7285 19907 7343 19913
rect 7285 19873 7297 19907
rect 7331 19904 7343 19907
rect 7466 19904 7472 19916
rect 7331 19876 7472 19904
rect 7331 19873 7343 19876
rect 7285 19867 7343 19873
rect 7466 19864 7472 19876
rect 7524 19864 7530 19916
rect 8202 19904 8208 19916
rect 8163 19876 8208 19904
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 8444 19876 9689 19904
rect 8444 19864 8450 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9950 19904 9956 19916
rect 9911 19876 9956 19904
rect 9677 19867 9735 19873
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 10410 19904 10416 19916
rect 10371 19876 10416 19904
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 10686 19904 10692 19916
rect 10647 19876 10692 19904
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 10796 19913 10824 20012
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 11977 20043 12035 20049
rect 11977 20040 11989 20043
rect 11388 20012 11989 20040
rect 11388 20000 11394 20012
rect 11977 20009 11989 20012
rect 12023 20009 12035 20043
rect 11977 20003 12035 20009
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13136 20012 13737 20040
rect 13136 20000 13142 20012
rect 13725 20009 13737 20012
rect 13771 20009 13783 20043
rect 13725 20003 13783 20009
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15436 20012 19012 20040
rect 15436 20000 15442 20012
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19873 10839 19907
rect 10781 19867 10839 19873
rect 6472 19808 7788 19836
rect 1946 19768 1952 19780
rect 1907 19740 1952 19768
rect 1946 19728 1952 19740
rect 2004 19728 2010 19780
rect 7760 19700 7788 19808
rect 7834 19796 7840 19848
rect 7892 19836 7898 19848
rect 11348 19836 11376 20000
rect 13354 19932 13360 19984
rect 13412 19972 13418 19984
rect 18322 19972 18328 19984
rect 13412 19944 14780 19972
rect 13412 19932 13418 19944
rect 11882 19904 11888 19916
rect 11843 19876 11888 19904
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19904 13139 19907
rect 13722 19904 13728 19916
rect 13127 19876 13728 19904
rect 13127 19873 13139 19876
rect 13081 19867 13139 19873
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 14752 19913 14780 19944
rect 16224 19944 18328 19972
rect 16224 19916 16252 19944
rect 18322 19932 18328 19944
rect 18380 19932 18386 19984
rect 18601 19975 18659 19981
rect 18601 19941 18613 19975
rect 18647 19972 18659 19975
rect 18690 19972 18696 19984
rect 18647 19944 18696 19972
rect 18647 19941 18659 19944
rect 18601 19935 18659 19941
rect 18690 19932 18696 19944
rect 18748 19932 18754 19984
rect 18984 19916 19012 20012
rect 21818 20000 21824 20052
rect 21876 20040 21882 20052
rect 22097 20043 22155 20049
rect 22097 20040 22109 20043
rect 21876 20012 22109 20040
rect 21876 20000 21882 20012
rect 22097 20009 22109 20012
rect 22143 20009 22155 20043
rect 22097 20003 22155 20009
rect 22646 20000 22652 20052
rect 22704 20040 22710 20052
rect 27062 20040 27068 20052
rect 22704 20012 27068 20040
rect 22704 20000 22710 20012
rect 27062 20000 27068 20012
rect 27120 20000 27126 20052
rect 20984 19975 21042 19981
rect 20984 19941 20996 19975
rect 21030 19972 21042 19975
rect 21174 19972 21180 19984
rect 21030 19944 21180 19972
rect 21030 19941 21042 19944
rect 20984 19935 21042 19941
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 22922 19932 22928 19984
rect 22980 19972 22986 19984
rect 23017 19975 23075 19981
rect 23017 19972 23029 19975
rect 22980 19944 23029 19972
rect 22980 19932 22986 19944
rect 23017 19941 23029 19944
rect 23063 19941 23075 19975
rect 23017 19935 23075 19941
rect 23566 19932 23572 19984
rect 23624 19972 23630 19984
rect 24118 19972 24124 19984
rect 23624 19944 24124 19972
rect 23624 19932 23630 19944
rect 24118 19932 24124 19944
rect 24176 19932 24182 19984
rect 14737 19907 14795 19913
rect 14737 19873 14749 19907
rect 14783 19873 14795 19907
rect 14737 19867 14795 19873
rect 15013 19907 15071 19913
rect 15013 19873 15025 19907
rect 15059 19904 15071 19907
rect 15286 19904 15292 19916
rect 15059 19876 15292 19904
rect 15059 19873 15071 19876
rect 15013 19867 15071 19873
rect 13446 19836 13452 19848
rect 7892 19808 11376 19836
rect 13407 19808 13452 19836
rect 7892 19796 7898 19808
rect 13446 19796 13452 19808
rect 13504 19836 13510 19848
rect 15028 19836 15056 19867
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 16206 19904 16212 19916
rect 16167 19876 16212 19904
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16476 19907 16534 19913
rect 16476 19873 16488 19907
rect 16522 19904 16534 19907
rect 17310 19904 17316 19916
rect 16522 19876 17316 19904
rect 16522 19873 16534 19876
rect 16476 19867 16534 19873
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 18414 19904 18420 19916
rect 18279 19876 18420 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 20073 19907 20131 19913
rect 20073 19904 20085 19907
rect 19024 19876 20085 19904
rect 19024 19864 19030 19876
rect 20073 19873 20085 19876
rect 20119 19873 20131 19907
rect 20073 19867 20131 19873
rect 22738 19864 22744 19916
rect 22796 19904 22802 19916
rect 22833 19907 22891 19913
rect 22833 19904 22845 19907
rect 22796 19876 22845 19904
rect 22796 19864 22802 19876
rect 22833 19873 22845 19876
rect 22879 19873 22891 19907
rect 22833 19867 22891 19873
rect 23109 19907 23167 19913
rect 23109 19873 23121 19907
rect 23155 19873 23167 19907
rect 23109 19867 23167 19873
rect 15470 19836 15476 19848
rect 13504 19808 15056 19836
rect 15431 19808 15476 19836
rect 13504 19796 13510 19808
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 19852 19808 20729 19836
rect 19852 19796 19858 19808
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 23124 19836 23152 19867
rect 23198 19864 23204 19916
rect 23256 19904 23262 19916
rect 23256 19876 23301 19904
rect 23256 19864 23262 19876
rect 23474 19864 23480 19916
rect 23532 19904 23538 19916
rect 23937 19907 23995 19913
rect 23937 19904 23949 19907
rect 23532 19876 23949 19904
rect 23532 19864 23538 19876
rect 23937 19873 23949 19876
rect 23983 19873 23995 19907
rect 23937 19867 23995 19873
rect 26044 19907 26102 19913
rect 26044 19873 26056 19907
rect 26090 19904 26102 19907
rect 26786 19904 26792 19916
rect 26090 19876 26792 19904
rect 26090 19873 26102 19876
rect 26044 19867 26102 19873
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 24578 19836 24584 19848
rect 23124 19808 24584 19836
rect 20717 19799 20775 19805
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 25774 19836 25780 19848
rect 25735 19808 25780 19836
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 10965 19771 11023 19777
rect 10965 19737 10977 19771
rect 11011 19768 11023 19771
rect 12710 19768 12716 19780
rect 11011 19740 12716 19768
rect 11011 19737 11023 19740
rect 10965 19731 11023 19737
rect 12710 19728 12716 19740
rect 12768 19728 12774 19780
rect 13262 19768 13268 19780
rect 13175 19740 13268 19768
rect 13261 19728 13268 19740
rect 13320 19768 13326 19780
rect 14090 19768 14096 19780
rect 13320 19740 14096 19768
rect 13320 19728 13326 19740
rect 14090 19728 14096 19740
rect 14148 19728 14154 19780
rect 14829 19771 14887 19777
rect 14829 19737 14841 19771
rect 14875 19768 14887 19771
rect 15010 19768 15016 19780
rect 14875 19740 15016 19768
rect 14875 19737 14887 19740
rect 14829 19731 14887 19737
rect 11054 19700 11060 19712
rect 7760 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 13078 19660 13084 19712
rect 13136 19700 13142 19712
rect 13261 19709 13289 19728
rect 13219 19703 13289 19709
rect 13219 19700 13231 19703
rect 13136 19672 13231 19700
rect 13136 19660 13142 19672
rect 13219 19669 13231 19672
rect 13265 19672 13289 19703
rect 13357 19703 13415 19709
rect 13265 19669 13277 19672
rect 13219 19663 13277 19669
rect 13357 19669 13369 19703
rect 13403 19700 13415 19703
rect 14844 19700 14872 19731
rect 15010 19728 15016 19740
rect 15068 19728 15074 19780
rect 20257 19771 20315 19777
rect 20257 19737 20269 19771
rect 20303 19768 20315 19771
rect 20346 19768 20352 19780
rect 20303 19740 20352 19768
rect 20303 19737 20315 19740
rect 20257 19731 20315 19737
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 17586 19700 17592 19712
rect 13403 19672 14872 19700
rect 17547 19672 17592 19700
rect 13403 19669 13415 19672
rect 13357 19663 13415 19669
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 23385 19703 23443 19709
rect 23385 19669 23397 19703
rect 23431 19700 23443 19703
rect 23566 19700 23572 19712
rect 23431 19672 23572 19700
rect 23431 19669 23443 19672
rect 23385 19663 23443 19669
rect 23566 19660 23572 19672
rect 23624 19660 23630 19712
rect 26694 19660 26700 19712
rect 26752 19700 26758 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 26752 19672 27169 19700
rect 26752 19660 26758 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 1104 19610 28428 19632
rect 1104 19558 5536 19610
rect 5588 19558 5600 19610
rect 5652 19558 5664 19610
rect 5716 19558 5728 19610
rect 5780 19558 14644 19610
rect 14696 19558 14708 19610
rect 14760 19558 14772 19610
rect 14824 19558 14836 19610
rect 14888 19558 23752 19610
rect 23804 19558 23816 19610
rect 23868 19558 23880 19610
rect 23932 19558 23944 19610
rect 23996 19558 28428 19610
rect 1104 19536 28428 19558
rect 2314 19456 2320 19508
rect 2372 19496 2378 19508
rect 9677 19499 9735 19505
rect 2372 19468 7604 19496
rect 2372 19456 2378 19468
rect 7576 19428 7604 19468
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 9950 19496 9956 19508
rect 9723 19468 9956 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 10413 19499 10471 19505
rect 10413 19465 10425 19499
rect 10459 19496 10471 19499
rect 10686 19496 10692 19508
rect 10459 19468 10692 19496
rect 10459 19465 10471 19468
rect 10413 19459 10471 19465
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 14001 19499 14059 19505
rect 14001 19496 14013 19499
rect 13780 19468 14013 19496
rect 13780 19456 13786 19468
rect 14001 19465 14013 19468
rect 14047 19465 14059 19499
rect 14001 19459 14059 19465
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19496 14427 19499
rect 14458 19496 14464 19508
rect 14415 19468 14464 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 17310 19496 17316 19508
rect 17271 19468 17316 19496
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 20441 19499 20499 19505
rect 17880 19468 20024 19496
rect 13078 19428 13084 19440
rect 7576 19400 13084 19428
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 13446 19388 13452 19440
rect 13504 19428 13510 19440
rect 13863 19431 13921 19437
rect 13863 19428 13875 19431
rect 13504 19400 13875 19428
rect 13504 19388 13510 19400
rect 13863 19397 13875 19400
rect 13909 19397 13921 19431
rect 15013 19431 15071 19437
rect 15013 19428 15025 19431
rect 13863 19391 13921 19397
rect 14016 19400 15025 19428
rect 10778 19360 10784 19372
rect 6656 19332 7144 19360
rect 1578 19252 1584 19304
rect 1636 19292 1642 19304
rect 3050 19292 3056 19304
rect 1636 19264 3056 19292
rect 1636 19252 1642 19264
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 5074 19292 5080 19304
rect 5035 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19292 5779 19295
rect 5902 19292 5908 19304
rect 5767 19264 5908 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 6270 19252 6276 19304
rect 6328 19292 6334 19304
rect 6454 19292 6460 19304
rect 6328 19264 6460 19292
rect 6328 19252 6334 19264
rect 6454 19252 6460 19264
rect 6512 19292 6518 19304
rect 6656 19292 6684 19332
rect 6822 19292 6828 19304
rect 6512 19264 6684 19292
rect 6783 19264 6828 19292
rect 6512 19252 6518 19264
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 7116 19301 7144 19332
rect 9508 19332 10784 19360
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 7101 19295 7159 19301
rect 7101 19261 7113 19295
rect 7147 19261 7159 19295
rect 7101 19255 7159 19261
rect 7193 19295 7251 19301
rect 7193 19261 7205 19295
rect 7239 19261 7251 19295
rect 7374 19292 7380 19304
rect 7335 19264 7380 19292
rect 7193 19255 7251 19261
rect 3320 19227 3378 19233
rect 3320 19193 3332 19227
rect 3366 19224 3378 19227
rect 4798 19224 4804 19236
rect 3366 19196 4804 19224
rect 3366 19193 3378 19196
rect 3320 19187 3378 19193
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 5169 19227 5227 19233
rect 5169 19193 5181 19227
rect 5215 19224 5227 19227
rect 7024 19224 7052 19255
rect 5215 19196 7052 19224
rect 7208 19224 7236 19255
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 8757 19295 8815 19301
rect 8757 19292 8769 19295
rect 7616 19264 8769 19292
rect 7616 19252 7622 19264
rect 8757 19261 8769 19264
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 9508 19292 9536 19332
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 11238 19360 11244 19372
rect 10980 19332 11244 19360
rect 8895 19264 9536 19292
rect 9585 19295 9643 19301
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9585 19261 9597 19295
rect 9631 19292 9643 19295
rect 9766 19292 9772 19304
rect 9631 19264 9772 19292
rect 9631 19261 9643 19264
rect 9585 19255 9643 19261
rect 9766 19252 9772 19264
rect 9824 19252 9830 19304
rect 10229 19295 10287 19301
rect 10229 19261 10241 19295
rect 10275 19292 10287 19295
rect 10980 19292 11008 19332
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 12805 19363 12863 19369
rect 12805 19329 12817 19363
rect 12851 19360 12863 19363
rect 12851 19332 13952 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 13924 19304 13952 19332
rect 11146 19292 11152 19304
rect 10275 19264 11008 19292
rect 11107 19264 11152 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 12250 19292 12256 19304
rect 11900 19264 12256 19292
rect 7834 19224 7840 19236
rect 7208 19196 7840 19224
rect 5215 19193 5227 19196
rect 5169 19187 5227 19193
rect 4433 19159 4491 19165
rect 4433 19125 4445 19159
rect 4479 19156 4491 19159
rect 4522 19156 4528 19168
rect 4479 19128 4528 19156
rect 4479 19125 4491 19128
rect 4433 19119 4491 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 5813 19159 5871 19165
rect 5813 19125 5825 19159
rect 5859 19156 5871 19159
rect 7006 19156 7012 19168
rect 5859 19128 7012 19156
rect 5859 19125 5871 19128
rect 5813 19119 5871 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7098 19116 7104 19168
rect 7156 19156 7162 19168
rect 7208 19156 7236 19196
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 11900 19224 11928 19264
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 13906 19252 13912 19304
rect 13964 19252 13970 19304
rect 10796 19196 11928 19224
rect 7156 19128 7236 19156
rect 7561 19159 7619 19165
rect 7156 19116 7162 19128
rect 7561 19125 7573 19159
rect 7607 19156 7619 19159
rect 8386 19156 8392 19168
rect 7607 19128 8392 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10796 19156 10824 19196
rect 11974 19184 11980 19236
rect 12032 19224 12038 19236
rect 12529 19227 12587 19233
rect 12529 19224 12541 19227
rect 12032 19196 12541 19224
rect 12032 19184 12038 19196
rect 12529 19193 12541 19196
rect 12575 19193 12587 19227
rect 12529 19187 12587 19193
rect 13725 19227 13783 19233
rect 13725 19193 13737 19227
rect 13771 19224 13783 19227
rect 14016 19224 14044 19400
rect 15013 19397 15025 19400
rect 15059 19428 15071 19431
rect 15746 19428 15752 19440
rect 15059 19400 15752 19428
rect 15059 19397 15071 19400
rect 15013 19391 15071 19397
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 17880 19428 17908 19468
rect 17644 19400 17908 19428
rect 19996 19428 20024 19468
rect 20441 19465 20453 19499
rect 20487 19496 20499 19499
rect 20714 19496 20720 19508
rect 20487 19468 20720 19496
rect 20487 19465 20499 19468
rect 20441 19459 20499 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 23198 19496 23204 19508
rect 22756 19468 23204 19496
rect 22646 19428 22652 19440
rect 19996 19400 22652 19428
rect 17644 19388 17650 19400
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 15102 19360 15108 19372
rect 14148 19332 15108 19360
rect 14148 19320 14154 19332
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 17788 19369 17816 19400
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 17773 19363 17831 19369
rect 17773 19329 17785 19363
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 17862 19320 17868 19372
rect 17920 19360 17926 19372
rect 17920 19332 17965 19360
rect 17920 19320 17926 19332
rect 20346 19320 20352 19372
rect 20404 19360 20410 19372
rect 20404 19332 21312 19360
rect 20404 19320 20410 19332
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 13771 19196 14044 19224
rect 14108 19264 14933 19292
rect 13771 19193 13783 19196
rect 13725 19187 13783 19193
rect 9732 19128 10824 19156
rect 9732 19116 9738 19128
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 10928 19128 10977 19156
rect 10928 19116 10934 19128
rect 10965 19125 10977 19128
rect 11011 19125 11023 19159
rect 10965 19119 11023 19125
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11606 19156 11612 19168
rect 11112 19128 11612 19156
rect 11112 19116 11118 19128
rect 11606 19116 11612 19128
rect 11664 19116 11670 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14108 19156 14136 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 15194 19292 15200 19304
rect 15155 19264 15200 19292
rect 14921 19255 14979 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 16117 19295 16175 19301
rect 16117 19292 16129 19295
rect 15804 19264 16129 19292
rect 15804 19252 15810 19264
rect 16117 19261 16129 19264
rect 16163 19261 16175 19295
rect 16117 19255 16175 19261
rect 18322 19252 18328 19304
rect 18380 19292 18386 19304
rect 18782 19292 18788 19304
rect 18380 19264 18788 19292
rect 18380 19252 18386 19264
rect 18782 19252 18788 19264
rect 18840 19292 18846 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18840 19264 19073 19292
rect 18840 19252 18846 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 20898 19292 20904 19304
rect 20680 19264 20904 19292
rect 20680 19252 20686 19264
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21284 19301 21312 19332
rect 21177 19295 21235 19301
rect 21177 19292 21189 19295
rect 21008 19264 21189 19292
rect 14734 19184 14740 19236
rect 14792 19224 14798 19236
rect 16209 19227 16267 19233
rect 16209 19224 16221 19227
rect 14792 19196 16221 19224
rect 14792 19184 14798 19196
rect 16209 19193 16221 19196
rect 16255 19193 16267 19227
rect 16209 19187 16267 19193
rect 19328 19227 19386 19233
rect 19328 19193 19340 19227
rect 19374 19224 19386 19227
rect 19374 19196 20576 19224
rect 19374 19193 19386 19196
rect 19328 19187 19386 19193
rect 13412 19128 14136 19156
rect 13412 19116 13418 19128
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 14516 19128 15393 19156
rect 14516 19116 14522 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 17126 19156 17132 19168
rect 17087 19128 17132 19156
rect 15381 19119 15439 19125
rect 17126 19116 17132 19128
rect 17184 19156 17190 19168
rect 17681 19159 17739 19165
rect 17681 19156 17693 19159
rect 17184 19128 17693 19156
rect 17184 19116 17190 19128
rect 17681 19125 17693 19128
rect 17727 19125 17739 19159
rect 20548 19156 20576 19196
rect 20714 19184 20720 19236
rect 20772 19224 20778 19236
rect 21008 19224 21036 19264
rect 21177 19261 21189 19264
rect 21223 19261 21235 19295
rect 21177 19255 21235 19261
rect 21269 19295 21327 19301
rect 21269 19261 21281 19295
rect 21315 19292 21327 19295
rect 22756 19292 22784 19468
rect 23198 19456 23204 19468
rect 23256 19456 23262 19508
rect 21315 19264 22784 19292
rect 22925 19295 22983 19301
rect 21315 19261 21327 19264
rect 21269 19255 21327 19261
rect 22925 19261 22937 19295
rect 22971 19292 22983 19295
rect 24765 19295 24823 19301
rect 24765 19292 24777 19295
rect 22971 19264 24777 19292
rect 22971 19261 22983 19264
rect 22925 19255 22983 19261
rect 24765 19261 24777 19264
rect 24811 19292 24823 19295
rect 25774 19292 25780 19304
rect 24811 19264 25780 19292
rect 24811 19261 24823 19264
rect 24765 19255 24823 19261
rect 20772 19196 21036 19224
rect 21085 19227 21143 19233
rect 20772 19184 20778 19196
rect 21085 19193 21097 19227
rect 21131 19224 21143 19227
rect 21358 19224 21364 19236
rect 21131 19196 21364 19224
rect 21131 19193 21143 19196
rect 21085 19187 21143 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 22554 19184 22560 19236
rect 22612 19224 22618 19236
rect 22940 19224 22968 19255
rect 25774 19252 25780 19264
rect 25832 19252 25838 19304
rect 26605 19295 26663 19301
rect 26605 19261 26617 19295
rect 26651 19292 26663 19295
rect 26694 19292 26700 19304
rect 26651 19264 26700 19292
rect 26651 19261 26663 19264
rect 26605 19255 26663 19261
rect 26694 19252 26700 19264
rect 26752 19292 26758 19304
rect 27338 19292 27344 19304
rect 26752 19264 27344 19292
rect 26752 19252 26758 19264
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 22612 19196 22968 19224
rect 23192 19227 23250 19233
rect 22612 19184 22618 19196
rect 23192 19193 23204 19227
rect 23238 19224 23250 19227
rect 23290 19224 23296 19236
rect 23238 19196 23296 19224
rect 23238 19193 23250 19196
rect 23192 19187 23250 19193
rect 23290 19184 23296 19196
rect 23348 19184 23354 19236
rect 23566 19184 23572 19236
rect 23624 19224 23630 19236
rect 25010 19227 25068 19233
rect 25010 19224 25022 19227
rect 23624 19196 25022 19224
rect 23624 19184 23630 19196
rect 25010 19193 25022 19196
rect 25056 19193 25068 19227
rect 25010 19187 25068 19193
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 20548 19128 21465 19156
rect 17681 19119 17739 19125
rect 21453 19125 21465 19128
rect 21499 19125 21511 19159
rect 21453 19119 21511 19125
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 22922 19156 22928 19168
rect 22520 19128 22928 19156
rect 22520 19116 22526 19128
rect 22922 19116 22928 19128
rect 22980 19116 22986 19168
rect 23014 19116 23020 19168
rect 23072 19156 23078 19168
rect 24305 19159 24363 19165
rect 24305 19156 24317 19159
rect 23072 19128 24317 19156
rect 23072 19116 23078 19128
rect 24305 19125 24317 19128
rect 24351 19156 24363 19159
rect 24486 19156 24492 19168
rect 24351 19128 24492 19156
rect 24351 19125 24363 19128
rect 24305 19119 24363 19125
rect 24486 19116 24492 19128
rect 24544 19116 24550 19168
rect 24578 19116 24584 19168
rect 24636 19156 24642 19168
rect 26145 19159 26203 19165
rect 26145 19156 26157 19159
rect 24636 19128 26157 19156
rect 24636 19116 24642 19128
rect 26145 19125 26157 19128
rect 26191 19125 26203 19159
rect 26145 19119 26203 19125
rect 1104 19066 28428 19088
rect 1104 19014 10090 19066
rect 10142 19014 10154 19066
rect 10206 19014 10218 19066
rect 10270 19014 10282 19066
rect 10334 19014 19198 19066
rect 19250 19014 19262 19066
rect 19314 19014 19326 19066
rect 19378 19014 19390 19066
rect 19442 19014 28428 19066
rect 1104 18992 28428 19014
rect 4798 18952 4804 18964
rect 4759 18924 4804 18952
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 6270 18912 6276 18964
rect 6328 18952 6334 18964
rect 7374 18952 7380 18964
rect 6328 18924 7380 18952
rect 6328 18912 6334 18924
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 9677 18955 9735 18961
rect 9677 18952 9689 18955
rect 7524 18924 9689 18952
rect 7524 18912 7530 18924
rect 9677 18921 9689 18924
rect 9723 18921 9735 18955
rect 14090 18952 14096 18964
rect 9677 18915 9735 18921
rect 13188 18924 14096 18952
rect 1489 18887 1547 18893
rect 1489 18853 1501 18887
rect 1535 18884 1547 18887
rect 2866 18884 2872 18896
rect 1535 18856 2872 18884
rect 1535 18853 1547 18856
rect 1489 18847 1547 18853
rect 2866 18844 2872 18856
rect 2924 18844 2930 18896
rect 4522 18884 4528 18896
rect 4483 18856 4528 18884
rect 4522 18844 4528 18856
rect 4580 18884 4586 18896
rect 5905 18887 5963 18893
rect 4580 18856 5304 18884
rect 4580 18844 4586 18856
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18816 2191 18819
rect 2314 18816 2320 18828
rect 2179 18788 2320 18816
rect 2179 18785 2191 18788
rect 2133 18779 2191 18785
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 4246 18816 4252 18828
rect 4207 18788 4252 18816
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 4430 18816 4436 18828
rect 4391 18788 4436 18816
rect 4430 18776 4436 18788
rect 4488 18776 4494 18828
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 4706 18816 4712 18828
rect 4663 18788 4712 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 5276 18825 5304 18856
rect 5905 18853 5917 18887
rect 5951 18884 5963 18887
rect 8941 18887 8999 18893
rect 5951 18856 8524 18884
rect 5951 18853 5963 18856
rect 5905 18847 5963 18853
rect 5261 18819 5319 18825
rect 5261 18785 5273 18819
rect 5307 18785 5319 18819
rect 5261 18779 5319 18785
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18816 6055 18819
rect 6086 18816 6092 18828
rect 6043 18788 6092 18816
rect 6043 18785 6055 18788
rect 5997 18779 6055 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18785 6239 18819
rect 6546 18816 6552 18828
rect 6507 18788 6552 18816
rect 6181 18779 6239 18785
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 6196 18748 6224 18779
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 6730 18776 6736 18828
rect 6788 18816 6794 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 6788 18788 7389 18816
rect 6788 18776 6794 18788
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 7377 18779 7435 18785
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18785 8079 18819
rect 8386 18816 8392 18828
rect 8347 18788 8392 18816
rect 8021 18779 8079 18785
rect 5399 18720 6224 18748
rect 6273 18751 6331 18757
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 6273 18717 6285 18751
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18748 6423 18751
rect 7098 18748 7104 18760
rect 6411 18720 7104 18748
rect 6411 18717 6423 18720
rect 6365 18711 6423 18717
rect 6288 18680 6316 18711
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 6454 18680 6460 18692
rect 6288 18652 6460 18680
rect 6454 18640 6460 18652
rect 6512 18640 6518 18692
rect 7193 18683 7251 18689
rect 7193 18680 7205 18683
rect 6564 18652 7205 18680
rect 1578 18612 1584 18624
rect 1539 18584 1584 18612
rect 1578 18572 1584 18584
rect 1636 18572 1642 18624
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 5905 18615 5963 18621
rect 5905 18612 5917 18615
rect 2556 18584 5917 18612
rect 2556 18572 2562 18584
rect 5905 18581 5917 18584
rect 5951 18581 5963 18615
rect 5905 18575 5963 18581
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6564 18612 6592 18652
rect 7193 18649 7205 18652
rect 7239 18649 7251 18683
rect 8036 18680 8064 18779
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8496 18816 8524 18856
rect 8941 18853 8953 18887
rect 8987 18884 8999 18887
rect 9585 18887 9643 18893
rect 9585 18884 9597 18887
rect 8987 18856 9597 18884
rect 8987 18853 8999 18856
rect 8941 18847 8999 18853
rect 9585 18853 9597 18856
rect 9631 18884 9643 18887
rect 12342 18884 12348 18896
rect 9631 18856 12348 18884
rect 9631 18853 9643 18856
rect 9585 18847 9643 18853
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 13188 18893 13216 18924
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18952 14243 18955
rect 18230 18952 18236 18964
rect 14231 18924 18236 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 20070 18912 20076 18964
rect 20128 18952 20134 18964
rect 23290 18952 23296 18964
rect 20128 18924 23152 18952
rect 23251 18924 23296 18952
rect 20128 18912 20134 18924
rect 13173 18887 13231 18893
rect 13173 18853 13185 18887
rect 13219 18853 13231 18887
rect 13173 18847 13231 18853
rect 13262 18844 13268 18896
rect 13320 18884 13326 18896
rect 17865 18887 17923 18893
rect 17865 18884 17877 18887
rect 13320 18856 17877 18884
rect 13320 18844 13326 18856
rect 17865 18853 17877 18856
rect 17911 18853 17923 18887
rect 17865 18847 17923 18853
rect 10226 18816 10232 18828
rect 8496 18788 10232 18816
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 10376 18788 10425 18816
rect 10376 18776 10382 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 11882 18816 11888 18828
rect 11843 18788 11888 18816
rect 10413 18779 10471 18785
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12986 18816 12992 18828
rect 12947 18788 12992 18816
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13354 18816 13360 18828
rect 13315 18788 13360 18816
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 14734 18816 14740 18828
rect 13964 18788 14740 18816
rect 13964 18776 13970 18788
rect 14734 18776 14740 18788
rect 14792 18776 14798 18828
rect 15010 18776 15016 18828
rect 15068 18816 15074 18828
rect 15930 18816 15936 18828
rect 15068 18788 15240 18816
rect 15891 18788 15936 18816
rect 15068 18776 15074 18788
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8343 18720 8953 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 8386 18680 8392 18692
rect 8036 18652 8392 18680
rect 7193 18643 7251 18649
rect 8386 18640 8392 18652
rect 8444 18640 8450 18692
rect 8481 18683 8539 18689
rect 8481 18649 8493 18683
rect 8527 18680 8539 18683
rect 9950 18680 9956 18692
rect 8527 18652 9956 18680
rect 8527 18649 8539 18652
rect 8481 18643 8539 18649
rect 9950 18640 9956 18652
rect 10008 18640 10014 18692
rect 10410 18640 10416 18692
rect 10468 18680 10474 18692
rect 10612 18680 10640 18711
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 14458 18748 14464 18760
rect 12308 18720 14464 18748
rect 12308 18708 12314 18720
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 15102 18748 15108 18760
rect 15063 18720 15108 18748
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15212 18748 15240 18788
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 16209 18819 16267 18825
rect 16209 18816 16221 18819
rect 16132 18788 16221 18816
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 15212 18720 16037 18748
rect 16025 18717 16037 18720
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 10468 18652 13676 18680
rect 10468 18640 10474 18652
rect 6144 18584 6592 18612
rect 6733 18615 6791 18621
rect 6144 18572 6150 18584
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 7098 18612 7104 18624
rect 6779 18584 7104 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 8113 18615 8171 18621
rect 8113 18612 8125 18615
rect 7432 18584 8125 18612
rect 7432 18572 7438 18584
rect 8113 18581 8125 18584
rect 8159 18581 8171 18615
rect 8113 18575 8171 18581
rect 9766 18572 9772 18624
rect 9824 18612 9830 18624
rect 10318 18612 10324 18624
rect 9824 18584 10324 18612
rect 9824 18572 9830 18584
rect 10318 18572 10324 18584
rect 10376 18612 10382 18624
rect 11974 18612 11980 18624
rect 10376 18584 11980 18612
rect 10376 18572 10382 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 13648 18612 13676 18652
rect 13722 18640 13728 18692
rect 13780 18680 13786 18692
rect 15013 18683 15071 18689
rect 15013 18680 15025 18683
rect 13780 18652 15025 18680
rect 13780 18640 13786 18652
rect 15013 18649 15025 18652
rect 15059 18649 15071 18683
rect 16132 18680 16160 18788
rect 16209 18785 16221 18788
rect 16255 18785 16267 18819
rect 16209 18779 16267 18785
rect 17129 18819 17187 18825
rect 17129 18785 17141 18819
rect 17175 18816 17187 18819
rect 17586 18816 17592 18828
rect 17175 18788 17592 18816
rect 17175 18785 17187 18788
rect 17129 18779 17187 18785
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 17770 18816 17776 18828
rect 17731 18788 17776 18816
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 18248 18825 18276 18912
rect 23014 18884 23020 18896
rect 18340 18856 22876 18884
rect 22975 18856 23020 18884
rect 18233 18819 18291 18825
rect 18233 18785 18245 18819
rect 18279 18785 18291 18819
rect 18233 18779 18291 18785
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18748 16543 18751
rect 17862 18748 17868 18760
rect 16531 18720 17868 18748
rect 16531 18717 16543 18720
rect 16485 18711 16543 18717
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 18340 18757 18368 18856
rect 18598 18816 18604 18828
rect 18559 18788 18604 18816
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 20070 18816 20076 18828
rect 18831 18788 20076 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 20248 18819 20306 18825
rect 20248 18785 20260 18819
rect 20294 18816 20306 18819
rect 20530 18816 20536 18828
rect 20294 18788 20536 18816
rect 20294 18785 20306 18788
rect 20248 18779 20306 18785
rect 20530 18776 20536 18788
rect 20588 18776 20594 18828
rect 20990 18776 20996 18828
rect 21048 18816 21054 18828
rect 22738 18816 22744 18828
rect 21048 18788 22744 18816
rect 21048 18776 21054 18788
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 19794 18708 19800 18760
rect 19852 18748 19858 18760
rect 19981 18751 20039 18757
rect 19981 18748 19993 18751
rect 19852 18720 19993 18748
rect 19852 18708 19858 18720
rect 19981 18717 19993 18720
rect 20027 18717 20039 18751
rect 22848 18748 22876 18856
rect 23014 18844 23020 18856
rect 23072 18844 23078 18896
rect 23124 18884 23152 18924
rect 23290 18912 23296 18924
rect 23348 18912 23354 18964
rect 24762 18912 24768 18964
rect 24820 18952 24826 18964
rect 26234 18952 26240 18964
rect 24820 18924 26240 18952
rect 24820 18912 24826 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 26786 18952 26792 18964
rect 26747 18924 26792 18952
rect 26786 18912 26792 18924
rect 26844 18912 26850 18964
rect 23124 18856 25268 18884
rect 22922 18776 22928 18828
rect 22980 18816 22986 18828
rect 23109 18819 23167 18825
rect 22980 18788 23025 18816
rect 22980 18776 22986 18788
rect 23109 18785 23121 18819
rect 23155 18816 23167 18819
rect 23198 18816 23204 18828
rect 23155 18788 23204 18816
rect 23155 18785 23167 18788
rect 23109 18779 23167 18785
rect 23198 18776 23204 18788
rect 23256 18776 23262 18828
rect 24121 18819 24179 18825
rect 24121 18785 24133 18819
rect 24167 18816 24179 18819
rect 24394 18816 24400 18828
rect 24167 18788 24400 18816
rect 24167 18785 24179 18788
rect 24121 18779 24179 18785
rect 24394 18776 24400 18788
rect 24452 18776 24458 18828
rect 25240 18825 25268 18856
rect 25314 18844 25320 18896
rect 25372 18884 25378 18896
rect 25501 18887 25559 18893
rect 25501 18884 25513 18887
rect 25372 18856 25513 18884
rect 25372 18844 25378 18856
rect 25501 18853 25513 18856
rect 25547 18853 25559 18887
rect 26970 18884 26976 18896
rect 25501 18847 25559 18853
rect 25608 18856 26976 18884
rect 25608 18825 25636 18856
rect 26970 18844 26976 18856
rect 27028 18844 27034 18896
rect 27522 18884 27528 18896
rect 27483 18856 27528 18884
rect 27522 18844 27528 18856
rect 27580 18844 27586 18896
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18785 25467 18819
rect 25409 18779 25467 18785
rect 25593 18819 25651 18825
rect 25593 18785 25605 18819
rect 25639 18785 25651 18819
rect 25593 18779 25651 18785
rect 24213 18751 24271 18757
rect 24213 18748 24225 18751
rect 22848 18720 24225 18748
rect 19981 18711 20039 18717
rect 24213 18717 24225 18720
rect 24259 18717 24271 18751
rect 24213 18711 24271 18717
rect 24486 18708 24492 18760
rect 24544 18748 24550 18760
rect 24762 18748 24768 18760
rect 24544 18720 24768 18748
rect 24544 18708 24550 18720
rect 24762 18708 24768 18720
rect 24820 18748 24826 18760
rect 25424 18748 25452 18779
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 26421 18819 26479 18825
rect 26292 18788 26337 18816
rect 26292 18776 26298 18788
rect 26421 18785 26433 18819
rect 26467 18785 26479 18819
rect 26421 18779 26479 18785
rect 26513 18819 26571 18825
rect 26513 18785 26525 18819
rect 26559 18785 26571 18819
rect 26513 18779 26571 18785
rect 26436 18748 26464 18779
rect 24820 18720 26464 18748
rect 24820 18708 24826 18720
rect 15013 18643 15071 18649
rect 15212 18652 16160 18680
rect 15212 18624 15240 18652
rect 24118 18640 24124 18692
rect 24176 18680 24182 18692
rect 26528 18680 26556 18779
rect 26602 18776 26608 18828
rect 26660 18816 26666 18828
rect 26660 18788 26705 18816
rect 26660 18776 26666 18788
rect 24176 18652 26556 18680
rect 24176 18640 24182 18652
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 13648 18584 14197 18612
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14185 18575 14243 18581
rect 14902 18615 14960 18621
rect 14902 18581 14914 18615
rect 14948 18612 14960 18615
rect 15194 18612 15200 18624
rect 14948 18584 15200 18612
rect 14948 18581 14960 18584
rect 14902 18575 14960 18581
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 15378 18612 15384 18624
rect 15339 18584 15384 18612
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 17221 18615 17279 18621
rect 17221 18612 17233 18615
rect 16632 18584 17233 18612
rect 16632 18572 16638 18584
rect 17221 18581 17233 18584
rect 17267 18581 17279 18615
rect 17221 18575 17279 18581
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 21361 18615 21419 18621
rect 21361 18612 21373 18615
rect 20312 18584 21373 18612
rect 20312 18572 20318 18584
rect 21361 18581 21373 18584
rect 21407 18581 21419 18615
rect 21361 18575 21419 18581
rect 25777 18615 25835 18621
rect 25777 18581 25789 18615
rect 25823 18612 25835 18615
rect 26234 18612 26240 18624
rect 25823 18584 26240 18612
rect 25823 18581 25835 18584
rect 25777 18575 25835 18581
rect 26234 18572 26240 18584
rect 26292 18572 26298 18624
rect 27614 18612 27620 18624
rect 27575 18584 27620 18612
rect 27614 18572 27620 18584
rect 27672 18572 27678 18624
rect 1104 18522 28428 18544
rect 1104 18470 5536 18522
rect 5588 18470 5600 18522
rect 5652 18470 5664 18522
rect 5716 18470 5728 18522
rect 5780 18470 14644 18522
rect 14696 18470 14708 18522
rect 14760 18470 14772 18522
rect 14824 18470 14836 18522
rect 14888 18470 23752 18522
rect 23804 18470 23816 18522
rect 23868 18470 23880 18522
rect 23932 18470 23944 18522
rect 23996 18470 28428 18522
rect 1104 18448 28428 18470
rect 4522 18408 4528 18420
rect 4435 18380 4528 18408
rect 4522 18368 4528 18380
rect 4580 18408 4586 18420
rect 5074 18408 5080 18420
rect 4580 18380 5080 18408
rect 4580 18368 4586 18380
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10686 18408 10692 18420
rect 9916 18380 10692 18408
rect 9916 18368 9922 18380
rect 10686 18368 10692 18380
rect 10744 18408 10750 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10744 18380 10977 18408
rect 10744 18368 10750 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 13173 18411 13231 18417
rect 13173 18377 13185 18411
rect 13219 18408 13231 18411
rect 13722 18408 13728 18420
rect 13219 18380 13728 18408
rect 13219 18377 13231 18380
rect 13173 18371 13231 18377
rect 13722 18368 13728 18380
rect 13780 18368 13786 18420
rect 18230 18408 18236 18420
rect 13832 18380 18236 18408
rect 6086 18340 6092 18352
rect 4448 18312 6092 18340
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 2866 18204 2872 18216
rect 2179 18176 2872 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 3050 18164 3056 18216
rect 3108 18204 3114 18216
rect 3145 18207 3203 18213
rect 3145 18204 3157 18207
rect 3108 18176 3157 18204
rect 3108 18164 3114 18176
rect 3145 18173 3157 18176
rect 3191 18204 3203 18207
rect 4448 18204 4476 18312
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 7561 18343 7619 18349
rect 7561 18309 7573 18343
rect 7607 18340 7619 18343
rect 7834 18340 7840 18352
rect 7607 18312 7840 18340
rect 7607 18309 7619 18312
rect 7561 18303 7619 18309
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 12986 18340 12992 18352
rect 10980 18312 12992 18340
rect 6362 18272 6368 18284
rect 5368 18244 6368 18272
rect 5368 18213 5396 18244
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 7006 18272 7012 18284
rect 6512 18244 6868 18272
rect 6967 18244 7012 18272
rect 6512 18232 6518 18244
rect 3191 18176 4476 18204
rect 5353 18207 5411 18213
rect 3191 18173 3203 18176
rect 3145 18167 3203 18173
rect 5353 18173 5365 18207
rect 5399 18173 5411 18207
rect 5353 18167 5411 18173
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18204 5779 18207
rect 5994 18204 6000 18216
rect 5767 18176 6000 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 5994 18164 6000 18176
rect 6052 18204 6058 18216
rect 6730 18204 6736 18216
rect 6052 18176 6736 18204
rect 6052 18164 6058 18176
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 6840 18204 6868 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 7374 18204 7380 18216
rect 6840 18176 7052 18204
rect 7335 18176 7380 18204
rect 1489 18139 1547 18145
rect 1489 18105 1501 18139
rect 1535 18136 1547 18139
rect 2038 18136 2044 18148
rect 1535 18108 2044 18136
rect 1535 18105 1547 18108
rect 1489 18099 1547 18105
rect 2038 18096 2044 18108
rect 2096 18096 2102 18148
rect 3412 18139 3470 18145
rect 3412 18105 3424 18139
rect 3458 18136 3470 18139
rect 4798 18136 4804 18148
rect 3458 18108 4804 18136
rect 3458 18105 3470 18108
rect 3412 18099 3470 18105
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 5537 18139 5595 18145
rect 5537 18105 5549 18139
rect 5583 18105 5595 18139
rect 5537 18099 5595 18105
rect 5629 18139 5687 18145
rect 5629 18105 5641 18139
rect 5675 18136 5687 18139
rect 6914 18136 6920 18148
rect 5675 18108 6920 18136
rect 5675 18105 5687 18108
rect 5629 18099 5687 18105
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 5552 18068 5580 18099
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 7024 18136 7052 18176
rect 7374 18164 7380 18176
rect 7432 18164 7438 18216
rect 7466 18164 7472 18216
rect 7524 18204 7530 18216
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 7524 18176 7573 18204
rect 7524 18164 7530 18176
rect 7561 18173 7573 18176
rect 7607 18173 7619 18207
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 7561 18167 7619 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18204 9643 18207
rect 10870 18204 10876 18216
rect 9631 18176 10876 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 9852 18139 9910 18145
rect 7024 18108 8432 18136
rect 5902 18068 5908 18080
rect 4672 18040 5580 18068
rect 5863 18040 5908 18068
rect 4672 18028 4678 18040
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 8404 18068 8432 18108
rect 9852 18105 9864 18139
rect 9898 18136 9910 18139
rect 10502 18136 10508 18148
rect 9898 18108 10508 18136
rect 9898 18105 9910 18108
rect 9852 18099 9910 18105
rect 10502 18096 10508 18108
rect 10560 18096 10566 18148
rect 10980 18068 11008 18312
rect 12986 18300 12992 18312
rect 13044 18340 13050 18352
rect 13044 18312 13124 18340
rect 13044 18300 13050 18312
rect 12084 18244 12664 18272
rect 12084 18213 12112 18244
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12250 18204 12256 18216
rect 12163 18176 12256 18204
rect 12069 18167 12127 18173
rect 11606 18096 11612 18148
rect 11664 18136 11670 18148
rect 12176 18136 12204 18176
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 12437 18207 12495 18213
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 12526 18204 12532 18216
rect 12483 18176 12532 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 12342 18136 12348 18148
rect 11664 18108 12204 18136
rect 12303 18108 12348 18136
rect 11664 18096 11670 18108
rect 12342 18096 12348 18108
rect 12400 18096 12406 18148
rect 12636 18136 12664 18244
rect 13096 18213 13124 18312
rect 13538 18300 13544 18352
rect 13596 18340 13602 18352
rect 13832 18340 13860 18380
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 19058 18408 19064 18420
rect 19019 18380 19064 18408
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 20530 18408 20536 18420
rect 20491 18380 20536 18408
rect 20530 18368 20536 18380
rect 20588 18368 20594 18420
rect 20990 18368 20996 18420
rect 21048 18408 21054 18420
rect 21177 18411 21235 18417
rect 21177 18408 21189 18411
rect 21048 18380 21189 18408
rect 21048 18368 21054 18380
rect 21177 18377 21189 18380
rect 21223 18377 21235 18411
rect 21177 18371 21235 18377
rect 24394 18368 24400 18420
rect 24452 18408 24458 18420
rect 27062 18408 27068 18420
rect 24452 18380 27068 18408
rect 24452 18368 24458 18380
rect 27062 18368 27068 18380
rect 27120 18368 27126 18420
rect 13596 18312 13860 18340
rect 14737 18343 14795 18349
rect 13596 18300 13602 18312
rect 14737 18309 14749 18343
rect 14783 18340 14795 18343
rect 15010 18340 15016 18352
rect 14783 18312 15016 18340
rect 14783 18309 14795 18312
rect 14737 18303 14795 18309
rect 15010 18300 15016 18312
rect 15068 18300 15074 18352
rect 15930 18300 15936 18352
rect 15988 18340 15994 18352
rect 18046 18340 18052 18352
rect 15988 18312 18052 18340
rect 15988 18300 15994 18312
rect 18046 18300 18052 18312
rect 18104 18340 18110 18352
rect 18104 18312 19334 18340
rect 18104 18300 18110 18312
rect 13354 18232 13360 18284
rect 13412 18232 13418 18284
rect 14458 18232 14464 18284
rect 14516 18272 14522 18284
rect 17957 18275 18015 18281
rect 17957 18272 17969 18275
rect 14516 18244 17969 18272
rect 14516 18232 14522 18244
rect 17957 18241 17969 18244
rect 18003 18272 18015 18275
rect 18598 18272 18604 18284
rect 18003 18244 18604 18272
rect 18003 18241 18015 18244
rect 17957 18235 18015 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 13081 18207 13139 18213
rect 13081 18173 13093 18207
rect 13127 18173 13139 18207
rect 13372 18204 13400 18232
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 13372 18176 14657 18204
rect 13081 18167 13139 18173
rect 14645 18173 14657 18176
rect 14691 18173 14703 18207
rect 14645 18167 14703 18173
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18204 14979 18207
rect 15102 18204 15108 18216
rect 14967 18176 15108 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15470 18164 15476 18216
rect 15528 18204 15534 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15528 18176 15853 18204
rect 15528 18164 15534 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 17773 18207 17831 18213
rect 17773 18173 17785 18207
rect 17819 18173 17831 18207
rect 17773 18167 17831 18173
rect 13262 18136 13268 18148
rect 12636 18108 13268 18136
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 13354 18096 13360 18148
rect 13412 18136 13418 18148
rect 13630 18136 13636 18148
rect 13412 18108 13636 18136
rect 13412 18096 13418 18108
rect 13630 18096 13636 18108
rect 13688 18136 13694 18148
rect 14001 18139 14059 18145
rect 14001 18136 14013 18139
rect 13688 18108 14013 18136
rect 13688 18096 13694 18108
rect 14001 18105 14013 18108
rect 14047 18105 14059 18139
rect 14001 18099 14059 18105
rect 15381 18139 15439 18145
rect 15381 18105 15393 18139
rect 15427 18136 15439 18139
rect 16758 18136 16764 18148
rect 15427 18108 16764 18136
rect 15427 18105 15439 18108
rect 15381 18099 15439 18105
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 17788 18136 17816 18167
rect 18414 18136 18420 18148
rect 17788 18108 18420 18136
rect 18414 18096 18420 18108
rect 18472 18136 18478 18148
rect 18785 18139 18843 18145
rect 18785 18136 18797 18139
rect 18472 18108 18797 18136
rect 18472 18096 18478 18108
rect 18785 18105 18797 18108
rect 18831 18105 18843 18139
rect 19306 18136 19334 18312
rect 19978 18300 19984 18352
rect 20036 18300 20042 18352
rect 22649 18343 22707 18349
rect 22649 18309 22661 18343
rect 22695 18340 22707 18343
rect 22695 18312 23980 18340
rect 22695 18309 22707 18312
rect 22649 18303 22707 18309
rect 19996 18272 20024 18300
rect 19996 18244 20162 18272
rect 19978 18204 19984 18216
rect 19939 18176 19984 18204
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20134 18213 20162 18244
rect 20119 18207 20177 18213
rect 20119 18173 20131 18207
rect 20165 18173 20177 18207
rect 20254 18204 20260 18216
rect 20215 18176 20260 18204
rect 20119 18167 20177 18173
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20404 18176 20449 18204
rect 20404 18164 20410 18176
rect 20622 18164 20628 18216
rect 20680 18204 20686 18216
rect 23952 18213 23980 18312
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18241 25467 18275
rect 25409 18235 25467 18241
rect 20993 18207 21051 18213
rect 20993 18204 21005 18207
rect 20680 18176 21005 18204
rect 20680 18164 20686 18176
rect 20993 18173 21005 18176
rect 21039 18173 21051 18207
rect 22833 18207 22891 18213
rect 22833 18204 22845 18207
rect 20993 18167 21051 18173
rect 22066 18176 22845 18204
rect 20530 18136 20536 18148
rect 19306 18108 20536 18136
rect 18785 18099 18843 18105
rect 20530 18096 20536 18108
rect 20588 18136 20594 18148
rect 22066 18136 22094 18176
rect 22833 18173 22845 18176
rect 22879 18173 22891 18207
rect 22833 18167 22891 18173
rect 23937 18207 23995 18213
rect 23937 18173 23949 18207
rect 23983 18204 23995 18207
rect 24302 18204 24308 18216
rect 23983 18176 24308 18204
rect 23983 18173 23995 18176
rect 23937 18167 23995 18173
rect 24302 18164 24308 18176
rect 24360 18164 24366 18216
rect 20588 18108 22094 18136
rect 20588 18096 20594 18108
rect 12618 18068 12624 18080
rect 8404 18040 11008 18068
rect 12579 18040 12624 18068
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 14093 18071 14151 18077
rect 14093 18037 14105 18071
rect 14139 18068 14151 18071
rect 14182 18068 14188 18080
rect 14139 18040 14188 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 16022 18068 16028 18080
rect 15935 18040 16028 18068
rect 16022 18028 16028 18040
rect 16080 18068 16086 18080
rect 16390 18068 16396 18080
rect 16080 18040 16396 18068
rect 16080 18028 16086 18040
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 17402 18028 17408 18080
rect 17460 18068 17466 18080
rect 21358 18068 21364 18080
rect 17460 18040 21364 18068
rect 17460 18028 17466 18040
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 22554 18028 22560 18080
rect 22612 18068 22618 18080
rect 23753 18071 23811 18077
rect 23753 18068 23765 18071
rect 22612 18040 23765 18068
rect 22612 18028 22618 18040
rect 23753 18037 23765 18040
rect 23799 18068 23811 18071
rect 25415 18068 25443 18235
rect 25590 18096 25596 18148
rect 25648 18145 25654 18148
rect 25648 18139 25712 18145
rect 25648 18105 25666 18139
rect 25700 18105 25712 18139
rect 25648 18099 25712 18105
rect 25648 18096 25654 18099
rect 25866 18068 25872 18080
rect 23799 18040 25872 18068
rect 23799 18037 23811 18040
rect 23753 18031 23811 18037
rect 25866 18028 25872 18040
rect 25924 18028 25930 18080
rect 26789 18071 26847 18077
rect 26789 18037 26801 18071
rect 26835 18068 26847 18071
rect 27338 18068 27344 18080
rect 26835 18040 27344 18068
rect 26835 18037 26847 18040
rect 26789 18031 26847 18037
rect 27338 18028 27344 18040
rect 27396 18028 27402 18080
rect 1104 17978 28428 18000
rect 1104 17926 10090 17978
rect 10142 17926 10154 17978
rect 10206 17926 10218 17978
rect 10270 17926 10282 17978
rect 10334 17926 19198 17978
rect 19250 17926 19262 17978
rect 19314 17926 19326 17978
rect 19378 17926 19390 17978
rect 19442 17926 28428 17978
rect 1104 17904 28428 17926
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 4798 17864 4804 17876
rect 3476 17836 4652 17864
rect 4759 17836 4804 17864
rect 3476 17824 3482 17836
rect 4522 17796 4528 17808
rect 4483 17768 4528 17796
rect 4522 17756 4528 17768
rect 4580 17756 4586 17808
rect 4624 17796 4652 17836
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 6972 17836 7113 17864
rect 6972 17824 6978 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 7101 17827 7159 17833
rect 4624 17768 4844 17796
rect 1848 17731 1906 17737
rect 1848 17697 1860 17731
rect 1894 17728 1906 17731
rect 4062 17728 4068 17740
rect 1894 17700 4068 17728
rect 1894 17697 1906 17700
rect 1848 17691 1906 17697
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4338 17737 4344 17740
rect 4295 17731 4344 17737
rect 4295 17697 4307 17731
rect 4341 17697 4344 17731
rect 4295 17691 4344 17697
rect 4338 17688 4344 17691
rect 4396 17688 4402 17740
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 4617 17731 4675 17737
rect 4617 17697 4629 17731
rect 4663 17728 4675 17731
rect 4706 17728 4712 17740
rect 4663 17700 4712 17728
rect 4663 17697 4675 17700
rect 4617 17691 4675 17697
rect 1394 17620 1400 17672
rect 1452 17660 1458 17672
rect 1581 17663 1639 17669
rect 1581 17660 1593 17663
rect 1452 17632 1593 17660
rect 1452 17620 1458 17632
rect 1581 17629 1593 17632
rect 1627 17629 1639 17663
rect 4448 17660 4476 17691
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 4816 17728 4844 17768
rect 5902 17756 5908 17808
rect 5960 17805 5966 17808
rect 5960 17799 6024 17805
rect 5960 17765 5978 17799
rect 6012 17765 6024 17799
rect 7116 17796 7144 17827
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7616 17836 7757 17864
rect 7616 17824 7622 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 8386 17864 8392 17876
rect 8347 17836 8392 17864
rect 7745 17827 7803 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 10502 17864 10508 17876
rect 10463 17836 10508 17864
rect 10502 17824 10508 17836
rect 10560 17824 10566 17876
rect 10962 17824 10968 17876
rect 11020 17864 11026 17876
rect 11020 17836 17264 17864
rect 11020 17824 11026 17836
rect 10137 17799 10195 17805
rect 7116 17768 8340 17796
rect 5960 17759 6024 17765
rect 5960 17756 5966 17759
rect 7653 17731 7711 17737
rect 4816 17700 6776 17728
rect 4522 17660 4528 17672
rect 4448 17632 4528 17660
rect 1581 17623 1639 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 1578 17484 1584 17536
rect 1636 17524 1642 17536
rect 2682 17524 2688 17536
rect 1636 17496 2688 17524
rect 1636 17484 1642 17496
rect 2682 17484 2688 17496
rect 2740 17524 2746 17536
rect 2961 17527 3019 17533
rect 2961 17524 2973 17527
rect 2740 17496 2973 17524
rect 2740 17484 2746 17496
rect 2961 17493 2973 17496
rect 3007 17493 3019 17527
rect 5736 17524 5764 17623
rect 6748 17592 6776 17700
rect 7653 17697 7665 17731
rect 7699 17728 7711 17731
rect 8202 17728 8208 17740
rect 7699 17700 8208 17728
rect 7699 17697 7711 17700
rect 7653 17691 7711 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 8312 17737 8340 17768
rect 10137 17765 10149 17799
rect 10183 17796 10195 17799
rect 11606 17796 11612 17808
rect 10183 17768 11612 17796
rect 10183 17765 10195 17768
rect 10137 17759 10195 17765
rect 11606 17756 11612 17768
rect 11664 17756 11670 17808
rect 11784 17799 11842 17805
rect 11784 17765 11796 17799
rect 11830 17796 11842 17799
rect 12618 17796 12624 17808
rect 11830 17768 12624 17796
rect 11830 17765 11842 17768
rect 11784 17759 11842 17765
rect 12618 17756 12624 17768
rect 12676 17756 12682 17808
rect 14366 17756 14372 17808
rect 14424 17796 14430 17808
rect 15013 17799 15071 17805
rect 15013 17796 15025 17799
rect 14424 17768 15025 17796
rect 14424 17756 14430 17768
rect 15013 17765 15025 17768
rect 15059 17765 15071 17799
rect 15013 17759 15071 17765
rect 16301 17799 16359 17805
rect 16301 17765 16313 17799
rect 16347 17796 16359 17799
rect 16482 17796 16488 17808
rect 16347 17768 16488 17796
rect 16347 17765 16359 17768
rect 16301 17759 16359 17765
rect 16482 17756 16488 17768
rect 16540 17756 16546 17808
rect 17236 17796 17264 17836
rect 18782 17824 18788 17876
rect 18840 17864 18846 17876
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 18840 17836 18889 17864
rect 18840 17824 18846 17836
rect 18877 17833 18889 17836
rect 18923 17833 18935 17867
rect 20070 17864 20076 17876
rect 20031 17836 20076 17864
rect 18877 17827 18935 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 26786 17864 26792 17876
rect 20824 17836 26792 17864
rect 20714 17796 20720 17808
rect 17236 17768 20720 17796
rect 20714 17756 20720 17768
rect 20772 17756 20778 17808
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17697 8355 17731
rect 9950 17728 9956 17740
rect 9911 17700 9956 17728
rect 8297 17691 8355 17697
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10229 17731 10287 17737
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17728 10379 17731
rect 10686 17728 10692 17740
rect 10367 17700 10692 17728
rect 10367 17697 10379 17700
rect 10321 17691 10379 17697
rect 10244 17660 10272 17691
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 10870 17688 10876 17740
rect 10928 17728 10934 17740
rect 11517 17731 11575 17737
rect 11517 17728 11529 17731
rect 10928 17700 11529 17728
rect 10928 17688 10934 17700
rect 11517 17697 11529 17700
rect 11563 17728 11575 17731
rect 12066 17728 12072 17740
rect 11563 17700 12072 17728
rect 11563 17697 11575 17700
rect 11517 17691 11575 17697
rect 12066 17688 12072 17700
rect 12124 17688 12130 17740
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17728 13691 17731
rect 13906 17728 13912 17740
rect 13679 17700 13912 17728
rect 13679 17697 13691 17700
rect 13633 17691 13691 17697
rect 13906 17688 13912 17700
rect 13964 17688 13970 17740
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14829 17731 14887 17737
rect 14829 17728 14841 17731
rect 14332 17700 14841 17728
rect 14332 17688 14338 17700
rect 14829 17697 14841 17700
rect 14875 17697 14887 17731
rect 14829 17691 14887 17697
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 15746 17728 15752 17740
rect 15611 17700 15752 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 16500 17728 16528 17756
rect 18598 17728 18604 17740
rect 16500 17700 18604 17728
rect 18598 17688 18604 17700
rect 18656 17688 18662 17740
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 19061 17731 19119 17737
rect 19061 17728 19073 17731
rect 18932 17700 19073 17728
rect 18932 17688 18938 17700
rect 19061 17697 19073 17700
rect 19107 17697 19119 17731
rect 19061 17691 19119 17697
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17728 20039 17731
rect 20254 17728 20260 17740
rect 20027 17700 20260 17728
rect 20027 17697 20039 17700
rect 19981 17691 20039 17697
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 10962 17660 10968 17672
rect 10244 17632 10968 17660
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 20824 17660 20852 17836
rect 26786 17824 26792 17836
rect 26844 17824 26850 17876
rect 22097 17799 22155 17805
rect 22097 17765 22109 17799
rect 22143 17796 22155 17799
rect 23474 17796 23480 17808
rect 22143 17768 23480 17796
rect 22143 17765 22155 17768
rect 22097 17759 22155 17765
rect 22112 17728 22140 17759
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 26234 17805 26240 17808
rect 26228 17796 26240 17805
rect 26195 17768 26240 17796
rect 26228 17759 26240 17768
rect 26234 17756 26240 17759
rect 26292 17756 26298 17808
rect 12676 17632 20852 17660
rect 21928 17700 22140 17728
rect 25317 17731 25375 17737
rect 12676 17620 12682 17632
rect 10870 17592 10876 17604
rect 6748 17564 10876 17592
rect 10870 17552 10876 17564
rect 10928 17552 10934 17604
rect 13817 17595 13875 17601
rect 12452 17564 13400 17592
rect 5994 17524 6000 17536
rect 5736 17496 6000 17524
rect 2961 17487 3019 17493
rect 5994 17484 6000 17496
rect 6052 17484 6058 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 12452 17524 12480 17564
rect 12308 17496 12480 17524
rect 12308 17484 12314 17496
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 12897 17527 12955 17533
rect 12897 17524 12909 17527
rect 12584 17496 12909 17524
rect 12584 17484 12590 17496
rect 12897 17493 12909 17496
rect 12943 17524 12955 17527
rect 13262 17524 13268 17536
rect 12943 17496 13268 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 13372 17524 13400 17564
rect 13817 17561 13829 17595
rect 13863 17592 13875 17595
rect 15010 17592 15016 17604
rect 13863 17564 15016 17592
rect 13863 17561 13875 17564
rect 13817 17555 13875 17561
rect 15010 17552 15016 17564
rect 15068 17552 15074 17604
rect 16485 17595 16543 17601
rect 16485 17592 16497 17595
rect 15120 17564 16497 17592
rect 14090 17524 14096 17536
rect 13372 17496 14096 17524
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 15120 17524 15148 17564
rect 16485 17561 16497 17564
rect 16531 17561 16543 17595
rect 16485 17555 16543 17561
rect 16666 17552 16672 17604
rect 16724 17592 16730 17604
rect 21928 17592 21956 17700
rect 25317 17697 25329 17731
rect 25363 17697 25375 17731
rect 25498 17728 25504 17740
rect 25459 17700 25504 17728
rect 25317 17691 25375 17697
rect 25332 17660 25360 17691
rect 25498 17688 25504 17700
rect 25556 17688 25562 17740
rect 25866 17688 25872 17740
rect 25924 17728 25930 17740
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 25924 17700 25973 17728
rect 25924 17688 25930 17700
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 25774 17660 25780 17672
rect 16724 17564 21956 17592
rect 22066 17632 25780 17660
rect 16724 17552 16730 17564
rect 14516 17496 15148 17524
rect 14516 17484 14522 17496
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15252 17496 15669 17524
rect 15252 17484 15258 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 18966 17524 18972 17536
rect 15804 17496 18972 17524
rect 15804 17484 15810 17496
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 22066 17524 22094 17632
rect 25774 17620 25780 17632
rect 25832 17620 25838 17672
rect 22186 17524 22192 17536
rect 19208 17496 22094 17524
rect 22147 17496 22192 17524
rect 19208 17484 19214 17496
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 26970 17484 26976 17536
rect 27028 17524 27034 17536
rect 27341 17527 27399 17533
rect 27341 17524 27353 17527
rect 27028 17496 27353 17524
rect 27028 17484 27034 17496
rect 27341 17493 27353 17496
rect 27387 17524 27399 17527
rect 27522 17524 27528 17536
rect 27387 17496 27528 17524
rect 27387 17493 27399 17496
rect 27341 17487 27399 17493
rect 27522 17484 27528 17496
rect 27580 17484 27586 17536
rect 1104 17434 28428 17456
rect 1104 17382 5536 17434
rect 5588 17382 5600 17434
rect 5652 17382 5664 17434
rect 5716 17382 5728 17434
rect 5780 17382 14644 17434
rect 14696 17382 14708 17434
rect 14760 17382 14772 17434
rect 14824 17382 14836 17434
rect 14888 17382 23752 17434
rect 23804 17382 23816 17434
rect 23868 17382 23880 17434
rect 23932 17382 23944 17434
rect 23996 17382 28428 17434
rect 1104 17360 28428 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 3050 17320 3056 17332
rect 1452 17292 3056 17320
rect 1452 17280 1458 17292
rect 1688 17193 1716 17292
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 4157 17323 4215 17329
rect 4157 17320 4169 17323
rect 4120 17292 4169 17320
rect 4120 17280 4126 17292
rect 4157 17289 4169 17292
rect 4203 17289 4215 17323
rect 4157 17283 4215 17289
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17320 4767 17323
rect 6546 17320 6552 17332
rect 4755 17292 6552 17320
rect 4755 17289 4767 17292
rect 4709 17283 4767 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 9122 17320 9128 17332
rect 6656 17292 9128 17320
rect 2774 17212 2780 17264
rect 2832 17252 2838 17264
rect 3970 17252 3976 17264
rect 2832 17224 3976 17252
rect 2832 17212 2838 17224
rect 3970 17212 3976 17224
rect 4028 17212 4034 17264
rect 4338 17212 4344 17264
rect 4396 17252 4402 17264
rect 5905 17255 5963 17261
rect 5905 17252 5917 17255
rect 4396 17224 5917 17252
rect 4396 17212 4402 17224
rect 5905 17221 5917 17224
rect 5951 17221 5963 17255
rect 5905 17215 5963 17221
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 6656 17184 6684 17292
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9858 17320 9864 17332
rect 9819 17292 9864 17320
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10594 17280 10600 17332
rect 10652 17320 10658 17332
rect 12526 17320 12532 17332
rect 10652 17292 12532 17320
rect 10652 17280 10658 17292
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 25590 17320 25596 17332
rect 15028 17292 19288 17320
rect 25551 17292 25596 17320
rect 7098 17252 7104 17264
rect 7059 17224 7104 17252
rect 7098 17212 7104 17224
rect 7156 17212 7162 17264
rect 7653 17255 7711 17261
rect 7653 17221 7665 17255
rect 7699 17252 7711 17255
rect 15028 17252 15056 17292
rect 7699 17224 15056 17252
rect 7699 17221 7711 17224
rect 7653 17215 7711 17221
rect 16206 17212 16212 17264
rect 16264 17252 16270 17264
rect 19150 17252 19156 17264
rect 16264 17224 19156 17252
rect 16264 17212 16270 17224
rect 19150 17212 19156 17224
rect 19208 17212 19214 17264
rect 8846 17184 8852 17196
rect 1673 17147 1731 17153
rect 3620 17156 6684 17184
rect 7208 17156 8852 17184
rect 3620 17128 3648 17156
rect 2682 17076 2688 17128
rect 2740 17116 2746 17128
rect 3602 17116 3608 17128
rect 2740 17088 3464 17116
rect 3515 17088 3608 17116
rect 2740 17076 2746 17088
rect 1940 17051 1998 17057
rect 1940 17017 1952 17051
rect 1986 17048 1998 17051
rect 3142 17048 3148 17060
rect 1986 17020 3148 17048
rect 1986 17017 1998 17020
rect 1940 17011 1998 17017
rect 3142 17008 3148 17020
rect 3200 17008 3206 17060
rect 3436 17048 3464 17088
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 3878 17116 3884 17128
rect 3712 17088 3884 17116
rect 3712 17048 3740 17088
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 4028 17088 4568 17116
rect 4028 17076 4034 17088
rect 3436 17020 3740 17048
rect 3789 17051 3847 17057
rect 3789 17017 3801 17051
rect 3835 17048 3847 17051
rect 4338 17048 4344 17060
rect 3835 17020 4344 17048
rect 3835 17017 3847 17020
rect 3789 17011 3847 17017
rect 4338 17008 4344 17020
rect 4396 17008 4402 17060
rect 4540 17048 4568 17088
rect 4614 17076 4620 17128
rect 4672 17116 4678 17128
rect 5721 17119 5779 17125
rect 4672 17088 4717 17116
rect 4672 17076 4678 17088
rect 5721 17085 5733 17119
rect 5767 17116 5779 17119
rect 7208 17116 7236 17156
rect 8846 17144 8852 17156
rect 8904 17184 8910 17196
rect 8904 17156 9996 17184
rect 8904 17144 8910 17156
rect 5767 17088 7236 17116
rect 7285 17119 7343 17125
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 7285 17085 7297 17119
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 7300 17048 7328 17079
rect 7374 17076 7380 17128
rect 7432 17116 7438 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7432 17088 7573 17116
rect 7432 17076 7438 17088
rect 7561 17085 7573 17088
rect 7607 17116 7619 17119
rect 8018 17116 8024 17128
rect 7607 17088 8024 17116
rect 7607 17085 7619 17088
rect 7561 17079 7619 17085
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 7466 17048 7472 17060
rect 4540 17020 4752 17048
rect 7300 17020 7472 17048
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3053 16983 3111 16989
rect 3053 16980 3065 16983
rect 3016 16952 3065 16980
rect 3016 16940 3022 16952
rect 3053 16949 3065 16952
rect 3099 16980 3111 16983
rect 4614 16980 4620 16992
rect 3099 16952 4620 16980
rect 3099 16949 3111 16952
rect 3053 16943 3111 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 4724 16980 4752 17020
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 7929 17051 7987 17057
rect 7929 17048 7941 17051
rect 7892 17020 7941 17048
rect 7892 17008 7898 17020
rect 7929 17017 7941 17020
rect 7975 17017 7987 17051
rect 9030 17048 9036 17060
rect 8991 17020 9036 17048
rect 7929 17011 7987 17017
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 9769 17051 9827 17057
rect 9769 17048 9781 17051
rect 9732 17020 9781 17048
rect 9732 17008 9738 17020
rect 9769 17017 9781 17020
rect 9815 17017 9827 17051
rect 9769 17011 9827 17017
rect 9858 16980 9864 16992
rect 4724 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 9968 16980 9996 17156
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12400 17156 15148 17184
rect 12400 17144 12406 17156
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 11940 17088 13553 17116
rect 11940 17076 11946 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 15120 17116 15148 17156
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 17678 17184 17684 17196
rect 17460 17156 17684 17184
rect 17460 17144 17466 17156
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17828 17156 17877 17184
rect 17828 17144 17834 17156
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 19260 17184 19288 17292
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 26878 17252 26884 17264
rect 20772 17224 25084 17252
rect 26839 17224 26884 17252
rect 20772 17212 20778 17224
rect 19610 17184 19616 17196
rect 19260 17156 19616 17184
rect 17865 17147 17923 17153
rect 19610 17144 19616 17156
rect 19668 17144 19674 17196
rect 22186 17184 22192 17196
rect 20640 17156 22192 17184
rect 20254 17116 20260 17128
rect 15120 17088 20260 17116
rect 15013 17079 15071 17085
rect 11514 17008 11520 17060
rect 11572 17048 11578 17060
rect 11572 17020 13860 17048
rect 11572 17008 11578 17020
rect 13538 16980 13544 16992
rect 9968 16952 13544 16980
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 13630 16940 13636 16992
rect 13688 16980 13694 16992
rect 13725 16983 13783 16989
rect 13725 16980 13737 16983
rect 13688 16952 13737 16980
rect 13688 16940 13694 16952
rect 13725 16949 13737 16952
rect 13771 16949 13783 16983
rect 13832 16980 13860 17020
rect 14182 17008 14188 17060
rect 14240 17048 14246 17060
rect 14369 17051 14427 17057
rect 14369 17048 14381 17051
rect 14240 17020 14381 17048
rect 14240 17008 14246 17020
rect 14369 17017 14381 17020
rect 14415 17017 14427 17051
rect 14369 17011 14427 17017
rect 14461 16983 14519 16989
rect 14461 16980 14473 16983
rect 13832 16952 14473 16980
rect 13725 16943 13783 16949
rect 14461 16949 14473 16952
rect 14507 16949 14519 16983
rect 15028 16980 15056 17079
rect 20254 17076 20260 17088
rect 20312 17076 20318 17128
rect 20640 17125 20668 17156
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 20349 17119 20407 17125
rect 20349 17085 20361 17119
rect 20395 17085 20407 17119
rect 20349 17079 20407 17085
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17085 20683 17119
rect 20625 17079 20683 17085
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17116 20775 17119
rect 21450 17116 21456 17128
rect 20763 17088 21456 17116
rect 20763 17085 20775 17088
rect 20717 17079 20775 17085
rect 15280 17051 15338 17057
rect 15280 17017 15292 17051
rect 15326 17048 15338 17051
rect 15470 17048 15476 17060
rect 15326 17020 15476 17048
rect 15326 17017 15338 17020
rect 15280 17011 15338 17017
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 16298 17008 16304 17060
rect 16356 17048 16362 17060
rect 16356 17020 17448 17048
rect 16356 17008 16362 17020
rect 17420 16992 17448 17020
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 20364 17048 20392 17079
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 21542 17076 21548 17128
rect 21600 17116 21606 17128
rect 22557 17119 22615 17125
rect 22557 17116 22569 17119
rect 21600 17088 22569 17116
rect 21600 17076 21606 17088
rect 22557 17085 22569 17088
rect 22603 17085 22615 17119
rect 22557 17079 22615 17085
rect 22925 17119 22983 17125
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 23934 17116 23940 17128
rect 22971 17088 23940 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 23934 17076 23940 17088
rect 23992 17076 23998 17128
rect 25056 17125 25084 17224
rect 26878 17212 26884 17224
rect 26936 17212 26942 17264
rect 27338 17184 27344 17196
rect 25424 17156 27344 17184
rect 25041 17119 25099 17125
rect 25041 17085 25053 17119
rect 25087 17085 25099 17119
rect 25314 17116 25320 17128
rect 25041 17079 25099 17085
rect 25148 17088 25320 17116
rect 18288 17020 20392 17048
rect 20533 17051 20591 17057
rect 18288 17008 18294 17020
rect 20533 17017 20545 17051
rect 20579 17048 20591 17051
rect 21082 17048 21088 17060
rect 20579 17020 21088 17048
rect 20579 17017 20591 17020
rect 20533 17011 20591 17017
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 22738 17048 22744 17060
rect 22699 17020 22744 17048
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 22833 17051 22891 17057
rect 22833 17017 22845 17051
rect 22879 17048 22891 17051
rect 25148 17048 25176 17088
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 25424 17125 25452 17156
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17085 25467 17119
rect 26694 17116 26700 17128
rect 26655 17088 26700 17116
rect 25409 17079 25467 17085
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 22879 17020 25176 17048
rect 25225 17051 25283 17057
rect 22879 17017 22891 17020
rect 22833 17011 22891 17017
rect 25225 17017 25237 17051
rect 25271 17017 25283 17051
rect 25225 17011 25283 17017
rect 15746 16980 15752 16992
rect 15028 16952 15752 16980
rect 14461 16943 14519 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 16393 16983 16451 16989
rect 16393 16949 16405 16983
rect 16439 16980 16451 16983
rect 16482 16980 16488 16992
rect 16439 16952 16488 16980
rect 16439 16949 16451 16952
rect 16393 16943 16451 16949
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 17310 16980 17316 16992
rect 17271 16952 17316 16980
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 17681 16983 17739 16989
rect 17681 16980 17693 16983
rect 17460 16952 17693 16980
rect 17460 16940 17466 16952
rect 17681 16949 17693 16952
rect 17727 16949 17739 16983
rect 17681 16943 17739 16949
rect 17773 16983 17831 16989
rect 17773 16949 17785 16983
rect 17819 16980 17831 16983
rect 17954 16980 17960 16992
rect 17819 16952 17960 16980
rect 17819 16949 17831 16952
rect 17773 16943 17831 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 20714 16980 20720 16992
rect 18104 16952 20720 16980
rect 18104 16940 18110 16952
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 20898 16980 20904 16992
rect 20859 16952 20904 16980
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 22848 16980 22876 17011
rect 23106 16980 23112 16992
rect 22520 16952 22876 16980
rect 23067 16952 23112 16980
rect 22520 16940 22526 16952
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 24946 16940 24952 16992
rect 25004 16980 25010 16992
rect 25240 16980 25268 17011
rect 25498 16980 25504 16992
rect 25004 16952 25504 16980
rect 25004 16940 25010 16952
rect 25498 16940 25504 16952
rect 25556 16940 25562 16992
rect 1104 16890 28428 16912
rect 1104 16838 10090 16890
rect 10142 16838 10154 16890
rect 10206 16838 10218 16890
rect 10270 16838 10282 16890
rect 10334 16838 19198 16890
rect 19250 16838 19262 16890
rect 19314 16838 19326 16890
rect 19378 16838 19390 16890
rect 19442 16838 28428 16890
rect 1104 16816 28428 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 1762 16776 1768 16788
rect 1627 16748 1768 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 2406 16736 2412 16788
rect 2464 16776 2470 16788
rect 3602 16776 3608 16788
rect 2464 16748 3608 16776
rect 2464 16736 2470 16748
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 2608 16640 2636 16748
rect 3602 16736 3608 16748
rect 3660 16736 3666 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 6270 16776 6276 16788
rect 4387 16748 6276 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 7834 16776 7840 16788
rect 7795 16748 7840 16776
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 10594 16776 10600 16788
rect 7944 16748 10600 16776
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 2958 16708 2964 16720
rect 2823 16680 2964 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 2958 16668 2964 16680
rect 3016 16668 3022 16720
rect 4430 16708 4436 16720
rect 3068 16680 4436 16708
rect 2547 16612 2636 16640
rect 2685 16643 2743 16649
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 2685 16609 2697 16643
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16609 2927 16643
rect 3068 16640 3096 16680
rect 4430 16668 4436 16680
rect 4488 16708 4494 16720
rect 5350 16708 5356 16720
rect 4488 16680 5356 16708
rect 4488 16668 4494 16680
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 6454 16708 6460 16720
rect 6052 16680 6460 16708
rect 6052 16668 6058 16680
rect 6454 16668 6460 16680
rect 6512 16668 6518 16720
rect 6638 16668 6644 16720
rect 6696 16708 6702 16720
rect 7944 16708 7972 16748
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 10870 16776 10876 16788
rect 10831 16748 10876 16776
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11020 16748 11529 16776
rect 11020 16736 11026 16748
rect 11517 16745 11529 16748
rect 11563 16776 11575 16779
rect 12342 16776 12348 16788
rect 11563 16748 12348 16776
rect 11563 16745 11575 16748
rect 11517 16739 11575 16745
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 15470 16776 15476 16788
rect 15335 16748 15476 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 16482 16776 16488 16788
rect 15948 16748 16488 16776
rect 12066 16708 12072 16720
rect 6696 16680 7972 16708
rect 9508 16680 12072 16708
rect 6696 16668 6702 16680
rect 2869 16603 2927 16609
rect 2976 16612 3096 16640
rect 2700 16504 2728 16603
rect 2774 16532 2780 16584
rect 2832 16572 2838 16584
rect 2884 16572 2912 16603
rect 2832 16544 2912 16572
rect 2832 16532 2838 16544
rect 2976 16504 3004 16612
rect 3142 16600 3148 16652
rect 3200 16600 3206 16652
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 3936 16612 4261 16640
rect 3936 16600 3942 16612
rect 4249 16609 4261 16612
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 2700 16476 3004 16504
rect 3053 16507 3111 16513
rect 3053 16473 3065 16507
rect 3099 16504 3111 16507
rect 3160 16504 3188 16600
rect 5912 16575 5970 16581
rect 5912 16541 5924 16575
rect 5958 16572 5970 16575
rect 6012 16572 6040 16668
rect 6172 16643 6230 16649
rect 6172 16609 6184 16643
rect 6218 16640 6230 16643
rect 7006 16640 7012 16652
rect 6218 16612 7012 16640
rect 6218 16609 6230 16612
rect 6172 16603 6230 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 9508 16649 9536 16680
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 12618 16708 12624 16720
rect 12579 16680 12624 16708
rect 12618 16668 12624 16680
rect 12676 16668 12682 16720
rect 12713 16711 12771 16717
rect 12713 16677 12725 16711
rect 12759 16708 12771 16711
rect 13446 16708 13452 16720
rect 12759 16680 13452 16708
rect 12759 16677 12771 16680
rect 12713 16671 12771 16677
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 15013 16711 15071 16717
rect 15013 16677 15025 16711
rect 15059 16708 15071 16711
rect 15948 16708 15976 16748
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17954 16776 17960 16788
rect 17175 16748 17960 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 18104 16748 18981 16776
rect 18104 16736 18110 16748
rect 18969 16745 18981 16748
rect 19015 16776 19027 16779
rect 19702 16776 19708 16788
rect 19015 16748 19708 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 21450 16736 21456 16788
rect 21508 16776 21514 16788
rect 21545 16779 21603 16785
rect 21545 16776 21557 16779
rect 21508 16748 21557 16776
rect 21508 16736 21514 16748
rect 21545 16745 21557 16748
rect 21591 16745 21603 16779
rect 23934 16776 23940 16788
rect 23847 16748 23940 16776
rect 21545 16739 21603 16745
rect 23934 16736 23940 16748
rect 23992 16776 23998 16788
rect 24486 16776 24492 16788
rect 23992 16748 24492 16776
rect 23992 16736 23998 16748
rect 24486 16736 24492 16748
rect 24544 16736 24550 16788
rect 25777 16779 25835 16785
rect 25777 16745 25789 16779
rect 25823 16776 25835 16779
rect 25866 16776 25872 16788
rect 25823 16748 25872 16776
rect 25823 16745 25835 16748
rect 25777 16739 25835 16745
rect 25866 16736 25872 16748
rect 25924 16736 25930 16788
rect 26142 16736 26148 16788
rect 26200 16776 26206 16788
rect 26421 16779 26479 16785
rect 26421 16776 26433 16779
rect 26200 16748 26433 16776
rect 26200 16736 26206 16748
rect 26421 16745 26433 16748
rect 26467 16745 26479 16779
rect 26421 16739 26479 16745
rect 15059 16680 15976 16708
rect 16016 16711 16074 16717
rect 15059 16677 15071 16680
rect 15013 16671 15071 16677
rect 16016 16677 16028 16711
rect 16062 16708 16074 16711
rect 17310 16708 17316 16720
rect 16062 16680 17316 16708
rect 16062 16677 16074 16680
rect 16016 16671 16074 16677
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 18782 16708 18788 16720
rect 17604 16680 18788 16708
rect 9766 16649 9772 16652
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16609 7803 16643
rect 7745 16603 7803 16609
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9760 16603 9772 16649
rect 9824 16640 9830 16652
rect 11425 16643 11483 16649
rect 9824 16612 9860 16640
rect 5958 16544 6040 16572
rect 5958 16541 5970 16544
rect 5912 16535 5970 16541
rect 3099 16476 3188 16504
rect 4264 16476 4476 16504
rect 3099 16473 3111 16476
rect 3053 16467 3111 16473
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 4264 16436 4292 16476
rect 1912 16408 4292 16436
rect 4448 16436 4476 16476
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 7285 16507 7343 16513
rect 7285 16504 7297 16507
rect 7156 16476 7297 16504
rect 7156 16464 7162 16476
rect 7285 16473 7297 16476
rect 7331 16504 7343 16507
rect 7760 16504 7788 16603
rect 9766 16600 9772 16603
rect 9824 16600 9830 16612
rect 11425 16609 11437 16643
rect 11471 16640 11483 16643
rect 11514 16640 11520 16652
rect 11471 16612 11520 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 12526 16640 12532 16652
rect 12483 16612 12532 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 12802 16640 12808 16652
rect 12763 16612 12808 16640
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 14458 16640 14464 16652
rect 13596 16612 14464 16640
rect 13596 16600 13602 16612
rect 14458 16600 14464 16612
rect 14516 16640 14522 16652
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14516 16612 14749 16640
rect 14516 16600 14522 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 15102 16640 15108 16652
rect 15063 16612 15108 16640
rect 14921 16603 14979 16609
rect 14936 16572 14964 16603
rect 15102 16600 15108 16612
rect 15160 16600 15166 16652
rect 15746 16640 15752 16652
rect 15659 16612 15752 16640
rect 15746 16600 15752 16612
rect 15804 16640 15810 16652
rect 17604 16649 17632 16680
rect 18782 16668 18788 16680
rect 18840 16668 18846 16720
rect 20432 16711 20490 16717
rect 20432 16677 20444 16711
rect 20478 16708 20490 16711
rect 20898 16708 20904 16720
rect 20478 16680 20904 16708
rect 20478 16677 20490 16680
rect 20432 16671 20490 16677
rect 20898 16668 20904 16680
rect 20956 16668 20962 16720
rect 22824 16711 22882 16717
rect 22824 16677 22836 16711
rect 22870 16708 22882 16711
rect 23106 16708 23112 16720
rect 22870 16680 23112 16708
rect 22870 16677 22882 16680
rect 22824 16671 22882 16677
rect 23106 16668 23112 16680
rect 23164 16668 23170 16720
rect 26329 16711 26387 16717
rect 26329 16677 26341 16711
rect 26375 16708 26387 16711
rect 26602 16708 26608 16720
rect 26375 16680 26608 16708
rect 26375 16677 26387 16680
rect 26329 16671 26387 16677
rect 26602 16668 26608 16680
rect 26660 16668 26666 16720
rect 17862 16649 17868 16652
rect 17589 16643 17647 16649
rect 17589 16640 17601 16643
rect 15804 16612 17601 16640
rect 15804 16600 15810 16612
rect 17589 16609 17601 16612
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 17856 16603 17868 16649
rect 17920 16640 17926 16652
rect 17920 16612 17956 16640
rect 17862 16600 17868 16603
rect 17920 16600 17926 16612
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 19852 16612 20177 16640
rect 19852 16600 19858 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 15010 16572 15016 16584
rect 14936 16544 15016 16572
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 7331 16476 7788 16504
rect 10428 16476 15792 16504
rect 7331 16473 7343 16476
rect 7285 16467 7343 16473
rect 10428 16436 10456 16476
rect 4448 16408 10456 16436
rect 1912 16396 1918 16408
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12768 16408 13001 16436
rect 12768 16396 12774 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 15764 16436 15792 16476
rect 20070 16436 20076 16448
rect 15764 16408 20076 16436
rect 12989 16399 13047 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20180 16436 20208 16603
rect 20254 16600 20260 16652
rect 20312 16640 20318 16652
rect 22462 16640 22468 16652
rect 20312 16612 22468 16640
rect 20312 16600 20318 16612
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 25590 16640 25596 16652
rect 25551 16612 25596 16640
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 25774 16600 25780 16652
rect 25832 16640 25838 16652
rect 26973 16643 27031 16649
rect 26973 16640 26985 16643
rect 25832 16612 26985 16640
rect 25832 16600 25838 16612
rect 26973 16609 26985 16612
rect 27019 16609 27031 16643
rect 26973 16603 27031 16609
rect 22554 16572 22560 16584
rect 22467 16544 22560 16572
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 22563 16436 22591 16532
rect 24578 16436 24584 16448
rect 20180 16408 24584 16436
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 1104 16346 28428 16368
rect 1104 16294 5536 16346
rect 5588 16294 5600 16346
rect 5652 16294 5664 16346
rect 5716 16294 5728 16346
rect 5780 16294 14644 16346
rect 14696 16294 14708 16346
rect 14760 16294 14772 16346
rect 14824 16294 14836 16346
rect 14888 16294 23752 16346
rect 23804 16294 23816 16346
rect 23868 16294 23880 16346
rect 23932 16294 23944 16346
rect 23996 16294 28428 16346
rect 1104 16272 28428 16294
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 15194 16232 15200 16244
rect 2188 16204 15200 16232
rect 2188 16192 2194 16204
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 18598 16192 18604 16244
rect 18656 16232 18662 16244
rect 18969 16235 19027 16241
rect 18969 16232 18981 16235
rect 18656 16204 18981 16232
rect 18656 16192 18662 16204
rect 18969 16201 18981 16204
rect 19015 16232 19027 16235
rect 20622 16232 20628 16244
rect 19015 16204 20628 16232
rect 19015 16201 19027 16204
rect 18969 16195 19027 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 21082 16192 21088 16244
rect 21140 16232 21146 16244
rect 21266 16232 21272 16244
rect 21140 16204 21272 16232
rect 21140 16192 21146 16204
rect 21266 16192 21272 16204
rect 21324 16232 21330 16244
rect 21545 16235 21603 16241
rect 21545 16232 21557 16235
rect 21324 16204 21557 16232
rect 21324 16192 21330 16204
rect 21545 16201 21557 16204
rect 21591 16201 21603 16235
rect 21545 16195 21603 16201
rect 22741 16235 22799 16241
rect 22741 16201 22753 16235
rect 22787 16232 22799 16235
rect 24762 16232 24768 16244
rect 22787 16204 24768 16232
rect 22787 16201 22799 16204
rect 22741 16195 22799 16201
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 25961 16235 26019 16241
rect 25961 16232 25973 16235
rect 25280 16204 25973 16232
rect 25280 16192 25286 16204
rect 25961 16201 25973 16204
rect 26007 16232 26019 16235
rect 26510 16232 26516 16244
rect 26007 16204 26516 16232
rect 26007 16201 26019 16204
rect 25961 16195 26019 16201
rect 26510 16192 26516 16204
rect 26568 16192 26574 16244
rect 5905 16167 5963 16173
rect 5905 16133 5917 16167
rect 5951 16164 5963 16167
rect 6362 16164 6368 16176
rect 5951 16136 6368 16164
rect 5951 16133 5963 16136
rect 5905 16127 5963 16133
rect 6362 16124 6368 16136
rect 6420 16124 6426 16176
rect 6454 16124 6460 16176
rect 6512 16164 6518 16176
rect 13446 16164 13452 16176
rect 6512 16136 8524 16164
rect 13407 16136 13452 16164
rect 6512 16124 6518 16136
rect 6086 16096 6092 16108
rect 3620 16068 6092 16096
rect 2038 15988 2044 16040
rect 2096 16028 2102 16040
rect 2133 16031 2191 16037
rect 2133 16028 2145 16031
rect 2096 16000 2145 16028
rect 2096 15988 2102 16000
rect 2133 15997 2145 16000
rect 2179 16028 2191 16031
rect 2222 16028 2228 16040
rect 2179 16000 2228 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 3620 16037 3648 16068
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 15997 3663 16031
rect 3786 16028 3792 16040
rect 3747 16000 3792 16028
rect 3605 15991 3663 15997
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 4632 16037 4660 16068
rect 6086 16056 6092 16068
rect 6144 16096 6150 16108
rect 6144 16068 6316 16096
rect 6144 16056 6150 16068
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 16028 4031 16031
rect 4617 16031 4675 16037
rect 4019 16000 4568 16028
rect 4019 15997 4031 16000
rect 3973 15991 4031 15997
rect 3881 15963 3939 15969
rect 3881 15929 3893 15963
rect 3927 15960 3939 15963
rect 4338 15960 4344 15972
rect 3927 15932 4344 15960
rect 3927 15929 3939 15932
rect 3881 15923 3939 15929
rect 4338 15920 4344 15932
rect 4396 15920 4402 15972
rect 4540 15960 4568 16000
rect 4617 15997 4629 16031
rect 4663 15997 4675 16031
rect 4985 16031 5043 16037
rect 4985 16028 4997 16031
rect 4617 15991 4675 15997
rect 4724 16000 4997 16028
rect 4724 15960 4752 16000
rect 4985 15997 4997 16000
rect 5031 16028 5043 16031
rect 5810 16028 5816 16040
rect 5031 16000 5816 16028
rect 5031 15997 5043 16000
rect 4985 15991 5043 15997
rect 5810 15988 5816 16000
rect 5868 15988 5874 16040
rect 4540 15932 4752 15960
rect 4801 15963 4859 15969
rect 4801 15929 4813 15963
rect 4847 15929 4859 15963
rect 4801 15923 4859 15929
rect 4154 15892 4160 15904
rect 4115 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 4816 15892 4844 15923
rect 4890 15920 4896 15972
rect 4948 15960 4954 15972
rect 5721 15963 5779 15969
rect 4948 15932 4993 15960
rect 4948 15920 4954 15932
rect 5721 15929 5733 15963
rect 5767 15960 5779 15963
rect 5902 15960 5908 15972
rect 5767 15932 5908 15960
rect 5767 15929 5779 15932
rect 5721 15923 5779 15929
rect 5902 15920 5908 15932
rect 5960 15920 5966 15972
rect 6288 15960 6316 16068
rect 6380 16028 6408 16124
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 8496 16105 8524 16136
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 15930 16164 15936 16176
rect 15891 16136 15936 16164
rect 15930 16124 15936 16136
rect 15988 16124 15994 16176
rect 16224 16136 17632 16164
rect 8481 16099 8539 16105
rect 6788 16068 7236 16096
rect 6788 16056 6794 16068
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6380 16000 6837 16028
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7098 16028 7104 16040
rect 7059 16000 7104 16028
rect 6825 15991 6883 15997
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 7208 16037 7236 16068
rect 8481 16065 8493 16099
rect 8527 16065 8539 16099
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 8481 16059 8539 16065
rect 13096 16068 14565 16096
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 15997 7251 16031
rect 12066 16028 12072 16040
rect 12027 16000 12072 16028
rect 7193 15991 7251 15997
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 12336 16031 12394 16037
rect 12336 15997 12348 16031
rect 12382 16028 12394 16031
rect 12710 16028 12716 16040
rect 12382 16000 12716 16028
rect 12382 15997 12394 16000
rect 12336 15991 12394 15997
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 13096 16028 13124 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 13004 16000 13124 16028
rect 6638 15960 6644 15972
rect 6288 15932 6644 15960
rect 6638 15920 6644 15932
rect 6696 15920 6702 15972
rect 7009 15963 7067 15969
rect 7009 15929 7021 15963
rect 7055 15960 7067 15963
rect 7834 15960 7840 15972
rect 7055 15932 7840 15960
rect 7055 15929 7067 15932
rect 7009 15923 7067 15929
rect 4982 15892 4988 15904
rect 4816 15864 4988 15892
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5350 15852 5356 15904
rect 5408 15892 5414 15904
rect 7024 15892 7052 15923
rect 7834 15920 7840 15932
rect 7892 15920 7898 15972
rect 8570 15920 8576 15972
rect 8628 15960 8634 15972
rect 8726 15963 8784 15969
rect 8726 15960 8738 15963
rect 8628 15932 8738 15960
rect 8628 15920 8634 15932
rect 8726 15929 8738 15932
rect 8772 15929 8784 15963
rect 8726 15923 8784 15929
rect 5408 15864 7052 15892
rect 5408 15852 5414 15864
rect 7098 15852 7104 15904
rect 7156 15892 7162 15904
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 7156 15864 7389 15892
rect 7156 15852 7162 15864
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 9858 15892 9864 15904
rect 9771 15864 9864 15892
rect 7377 15855 7435 15861
rect 9858 15852 9864 15864
rect 9916 15892 9922 15904
rect 13004 15892 13032 16000
rect 13446 15988 13452 16040
rect 13504 16028 13510 16040
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 13504 16000 13921 16028
rect 13504 15988 13510 16000
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 16028 14703 16031
rect 16224 16028 16252 16136
rect 17604 16096 17632 16136
rect 17862 16124 17868 16176
rect 17920 16164 17926 16176
rect 17920 16136 17965 16164
rect 17920 16124 17926 16136
rect 18230 16124 18236 16176
rect 18288 16164 18294 16176
rect 23382 16164 23388 16176
rect 18288 16136 23388 16164
rect 18288 16124 18294 16136
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 24578 16096 24584 16108
rect 17604 16068 23612 16096
rect 24539 16068 24584 16096
rect 14691 16000 16252 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 17313 16031 17371 16037
rect 17313 16028 17325 16031
rect 16356 16000 17325 16028
rect 16356 15988 16362 16000
rect 17313 15997 17325 16000
rect 17359 15997 17371 16031
rect 17313 15991 17371 15997
rect 17681 16031 17739 16037
rect 17681 15997 17693 16031
rect 17727 16028 17739 16031
rect 17862 16028 17868 16040
rect 17727 16000 17868 16028
rect 17727 15997 17739 16000
rect 17681 15991 17739 15997
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18656 16000 18889 16028
rect 18656 15988 18662 16000
rect 18877 15997 18889 16000
rect 18923 16028 18935 16031
rect 18966 16028 18972 16040
rect 18923 16000 18972 16028
rect 18923 15997 18935 16000
rect 18877 15991 18935 15997
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 19521 16031 19579 16037
rect 19521 15997 19533 16031
rect 19567 15997 19579 16031
rect 19521 15991 19579 15997
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 17402 15960 17408 15972
rect 15068 15932 17408 15960
rect 15068 15920 15074 15932
rect 17402 15920 17408 15932
rect 17460 15960 17466 15972
rect 17497 15963 17555 15969
rect 17497 15960 17509 15963
rect 17460 15932 17509 15960
rect 17460 15920 17466 15932
rect 17497 15929 17509 15932
rect 17543 15929 17555 15963
rect 17497 15923 17555 15929
rect 17589 15963 17647 15969
rect 17589 15929 17601 15963
rect 17635 15960 17647 15963
rect 18046 15960 18052 15972
rect 17635 15932 18052 15960
rect 17635 15929 17647 15932
rect 17589 15923 17647 15929
rect 18046 15920 18052 15932
rect 18104 15960 18110 15972
rect 18322 15960 18328 15972
rect 18104 15932 18328 15960
rect 18104 15920 18110 15932
rect 18322 15920 18328 15932
rect 18380 15920 18386 15972
rect 19536 15960 19564 15991
rect 19610 15988 19616 16040
rect 19668 16028 19674 16040
rect 20438 16028 20444 16040
rect 19668 16000 20444 16028
rect 19668 15988 19674 16000
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 16028 23443 16031
rect 23474 16028 23480 16040
rect 23431 16000 23480 16028
rect 23431 15997 23443 16000
rect 23385 15991 23443 15997
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 23584 16028 23612 16068
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 25314 16028 25320 16040
rect 23584 16000 25320 16028
rect 25314 15988 25320 16000
rect 25372 15988 25378 16040
rect 19702 15960 19708 15972
rect 19536 15932 19708 15960
rect 19702 15920 19708 15932
rect 19760 15960 19766 15972
rect 20898 15960 20904 15972
rect 19760 15932 20904 15960
rect 19760 15920 19766 15932
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 20990 15920 20996 15972
rect 21048 15960 21054 15972
rect 21453 15963 21511 15969
rect 21453 15960 21465 15963
rect 21048 15932 21465 15960
rect 21048 15920 21054 15932
rect 21453 15929 21465 15932
rect 21499 15960 21511 15963
rect 21910 15960 21916 15972
rect 21499 15932 21916 15960
rect 21499 15929 21511 15932
rect 21453 15923 21511 15929
rect 21910 15920 21916 15932
rect 21968 15960 21974 15972
rect 22649 15963 22707 15969
rect 22649 15960 22661 15963
rect 21968 15932 22661 15960
rect 21968 15920 21974 15932
rect 22649 15929 22661 15932
rect 22695 15929 22707 15963
rect 23566 15960 23572 15972
rect 23527 15932 23572 15960
rect 22649 15923 22707 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 24854 15969 24860 15972
rect 24848 15923 24860 15969
rect 24912 15960 24918 15972
rect 26697 15963 26755 15969
rect 24912 15932 24948 15960
rect 24854 15920 24860 15923
rect 24912 15920 24918 15932
rect 26697 15929 26709 15963
rect 26743 15960 26755 15963
rect 26878 15960 26884 15972
rect 26743 15932 26884 15960
rect 26743 15929 26755 15932
rect 26697 15923 26755 15929
rect 26878 15920 26884 15932
rect 26936 15920 26942 15972
rect 9916 15864 13032 15892
rect 9916 15852 9922 15864
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14001 15895 14059 15901
rect 14001 15892 14013 15895
rect 13780 15864 14013 15892
rect 13780 15852 13786 15864
rect 14001 15861 14013 15864
rect 14047 15861 14059 15895
rect 14001 15855 14059 15861
rect 14553 15895 14611 15901
rect 14553 15861 14565 15895
rect 14599 15892 14611 15895
rect 20806 15892 20812 15904
rect 14599 15864 20812 15892
rect 14599 15861 14611 15864
rect 14553 15855 14611 15861
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 22278 15852 22284 15904
rect 22336 15892 22342 15904
rect 26789 15895 26847 15901
rect 26789 15892 26801 15895
rect 22336 15864 26801 15892
rect 22336 15852 22342 15864
rect 26789 15861 26801 15864
rect 26835 15861 26847 15895
rect 26789 15855 26847 15861
rect 1104 15802 28428 15824
rect 1104 15750 10090 15802
rect 10142 15750 10154 15802
rect 10206 15750 10218 15802
rect 10270 15750 10282 15802
rect 10334 15750 19198 15802
rect 19250 15750 19262 15802
rect 19314 15750 19326 15802
rect 19378 15750 19390 15802
rect 19442 15750 28428 15802
rect 1104 15728 28428 15750
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 5994 15688 6000 15700
rect 2372 15660 6000 15688
rect 2372 15648 2378 15660
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 6328 15660 9536 15688
rect 6328 15648 6334 15660
rect 4516 15623 4574 15629
rect 4516 15589 4528 15623
rect 4562 15620 4574 15623
rect 5166 15620 5172 15632
rect 4562 15592 5172 15620
rect 4562 15589 4574 15592
rect 4516 15583 4574 15589
rect 5166 15580 5172 15592
rect 5224 15580 5230 15632
rect 6730 15580 6736 15632
rect 6788 15620 6794 15632
rect 6825 15623 6883 15629
rect 6825 15620 6837 15623
rect 6788 15592 6837 15620
rect 6788 15580 6794 15592
rect 6825 15589 6837 15592
rect 6871 15589 6883 15623
rect 6825 15583 6883 15589
rect 7282 15580 7288 15632
rect 7340 15620 7346 15632
rect 7377 15623 7435 15629
rect 7377 15620 7389 15623
rect 7340 15592 7389 15620
rect 7340 15580 7346 15592
rect 7377 15589 7389 15592
rect 7423 15589 7435 15623
rect 7377 15583 7435 15589
rect 7650 15580 7656 15632
rect 7708 15620 7714 15632
rect 8573 15623 8631 15629
rect 8573 15620 8585 15623
rect 7708 15592 8585 15620
rect 7708 15580 7714 15592
rect 8573 15589 8585 15592
rect 8619 15589 8631 15623
rect 8573 15583 8631 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15552 4307 15555
rect 6454 15552 6460 15564
rect 4295 15524 6460 15552
rect 4295 15521 4307 15524
rect 4249 15515 4307 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 6914 15552 6920 15564
rect 6687 15524 6920 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 9508 15561 9536 15660
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 9824 15660 10057 15688
rect 9824 15648 9830 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10744 15660 22094 15688
rect 10744 15648 10750 15660
rect 9677 15623 9735 15629
rect 9677 15589 9689 15623
rect 9723 15620 9735 15623
rect 12894 15620 12900 15632
rect 9723 15592 12900 15620
rect 9723 15589 9735 15592
rect 9677 15583 9735 15589
rect 12894 15580 12900 15592
rect 12952 15580 12958 15632
rect 14366 15620 14372 15632
rect 13464 15592 14372 15620
rect 10870 15561 10876 15564
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15521 9551 15555
rect 9493 15515 9551 15521
rect 9769 15555 9827 15561
rect 9769 15521 9781 15555
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15552 9919 15555
rect 10856 15555 10876 15561
rect 9907 15524 10824 15552
rect 9907 15521 9919 15524
rect 9861 15515 9919 15521
rect 5810 15376 5816 15428
rect 5868 15416 5874 15428
rect 8404 15416 8432 15515
rect 9784 15484 9812 15515
rect 10686 15484 10692 15496
rect 9784 15456 10692 15484
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 10796 15484 10824 15524
rect 10856 15521 10868 15555
rect 10856 15515 10876 15521
rect 10870 15512 10876 15515
rect 10928 15512 10934 15564
rect 13354 15552 13360 15564
rect 13315 15524 13360 15552
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 13464 15561 13492 15592
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 16482 15580 16488 15632
rect 16540 15620 16546 15632
rect 16540 15592 18828 15620
rect 16540 15580 16546 15592
rect 13449 15555 13507 15561
rect 13449 15521 13461 15555
rect 13495 15521 13507 15555
rect 13722 15552 13728 15564
rect 13683 15524 13728 15552
rect 13449 15515 13507 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 15004 15555 15062 15561
rect 15004 15521 15016 15555
rect 15050 15552 15062 15555
rect 15286 15552 15292 15564
rect 15050 15524 15292 15552
rect 15050 15521 15062 15524
rect 15004 15515 15062 15521
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 17034 15552 17040 15564
rect 16899 15524 17040 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 17034 15512 17040 15524
rect 17092 15512 17098 15564
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15521 17555 15555
rect 17497 15515 17555 15521
rect 10962 15484 10968 15496
rect 10796 15456 10968 15484
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 12066 15444 12072 15496
rect 12124 15484 12130 15496
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 12124 15456 14749 15484
rect 12124 15444 12130 15456
rect 14737 15453 14749 15456
rect 14783 15453 14795 15487
rect 17512 15484 17540 15515
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18800 15561 18828 15592
rect 20070 15580 20076 15632
rect 20128 15620 20134 15632
rect 21910 15620 21916 15632
rect 20128 15592 20484 15620
rect 21871 15592 21916 15620
rect 20128 15580 20134 15592
rect 20254 15561 20260 15564
rect 18141 15555 18199 15561
rect 18141 15552 18153 15555
rect 18012 15524 18153 15552
rect 18012 15512 18018 15524
rect 18141 15521 18153 15524
rect 18187 15521 18199 15555
rect 18141 15515 18199 15521
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 20248 15515 20260 15561
rect 20312 15552 20318 15564
rect 20456 15552 20484 15592
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 22066 15620 22094 15660
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23937 15691 23995 15697
rect 23937 15688 23949 15691
rect 23440 15660 23949 15688
rect 23440 15648 23446 15660
rect 23937 15657 23949 15660
rect 23983 15657 23995 15691
rect 23937 15651 23995 15657
rect 26510 15648 26516 15700
rect 26568 15688 26574 15700
rect 26605 15691 26663 15697
rect 26605 15688 26617 15691
rect 26568 15660 26617 15688
rect 26568 15648 26574 15660
rect 26605 15657 26617 15660
rect 26651 15688 26663 15691
rect 27246 15688 27252 15700
rect 26651 15660 27252 15688
rect 26651 15657 26663 15660
rect 26605 15651 26663 15657
rect 27246 15648 27252 15660
rect 27304 15648 27310 15700
rect 25590 15620 25596 15632
rect 22066 15592 25596 15620
rect 25590 15580 25596 15592
rect 25648 15620 25654 15632
rect 27341 15623 27399 15629
rect 27341 15620 27353 15623
rect 25648 15592 27353 15620
rect 25648 15580 25654 15592
rect 27341 15589 27353 15592
rect 27387 15589 27399 15623
rect 27341 15583 27399 15589
rect 22824 15555 22882 15561
rect 20312 15524 20348 15552
rect 20456 15524 21404 15552
rect 20254 15512 20260 15515
rect 20312 15512 20318 15524
rect 14737 15447 14795 15453
rect 16132 15456 17540 15484
rect 19981 15487 20039 15493
rect 9030 15416 9036 15428
rect 5868 15388 7512 15416
rect 8404 15388 9036 15416
rect 5868 15376 5874 15388
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 2314 15348 2320 15360
rect 1627 15320 2320 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 4890 15308 4896 15360
rect 4948 15348 4954 15360
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 4948 15320 5641 15348
rect 4948 15308 4954 15320
rect 5629 15317 5641 15320
rect 5675 15348 5687 15351
rect 6178 15348 6184 15360
rect 5675 15320 6184 15348
rect 5675 15317 5687 15320
rect 5629 15311 5687 15317
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 7484 15357 7512 15388
rect 9030 15376 9036 15388
rect 9088 15416 9094 15428
rect 10870 15416 10876 15428
rect 9088 15388 10876 15416
rect 9088 15376 9094 15388
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 11054 15416 11060 15428
rect 11015 15388 11060 15416
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 14182 15376 14188 15428
rect 14240 15416 14246 15428
rect 14240 15388 14596 15416
rect 14240 15376 14246 15388
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 12802 15348 12808 15360
rect 7515 15320 12808 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13170 15348 13176 15360
rect 13131 15320 13176 15348
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13633 15351 13691 15357
rect 13633 15317 13645 15351
rect 13679 15348 13691 15351
rect 13814 15348 13820 15360
rect 13679 15320 13820 15348
rect 13679 15317 13691 15320
rect 13633 15311 13691 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14568 15348 14596 15388
rect 15746 15376 15752 15428
rect 15804 15416 15810 15428
rect 16132 15425 16160 15456
rect 19981 15453 19993 15487
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 16117 15419 16175 15425
rect 16117 15416 16129 15419
rect 15804 15388 16129 15416
rect 15804 15376 15810 15388
rect 16117 15385 16129 15388
rect 16163 15385 16175 15419
rect 17218 15416 17224 15428
rect 16117 15379 16175 15385
rect 16960 15388 17224 15416
rect 16960 15357 16988 15388
rect 17218 15376 17224 15388
rect 17276 15416 17282 15428
rect 17862 15416 17868 15428
rect 17276 15388 17868 15416
rect 17276 15376 17282 15388
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 16945 15351 17003 15357
rect 16945 15348 16957 15351
rect 14568 15320 16957 15348
rect 16945 15317 16957 15320
rect 16991 15317 17003 15351
rect 16945 15311 17003 15317
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 17589 15351 17647 15357
rect 17589 15348 17601 15351
rect 17460 15320 17601 15348
rect 17460 15308 17466 15320
rect 17589 15317 17601 15320
rect 17635 15317 17647 15351
rect 17589 15311 17647 15317
rect 18046 15308 18052 15360
rect 18104 15348 18110 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18104 15320 18245 15348
rect 18104 15308 18110 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18874 15348 18880 15360
rect 18835 15320 18880 15348
rect 18233 15311 18291 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19996 15348 20024 15447
rect 21376 15425 21404 15524
rect 22824 15521 22836 15555
rect 22870 15552 22882 15555
rect 23382 15552 23388 15564
rect 22870 15524 23388 15552
rect 22870 15521 22882 15524
rect 22824 15515 22882 15521
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 24946 15512 24952 15564
rect 25004 15552 25010 15564
rect 25481 15555 25539 15561
rect 25481 15552 25493 15555
rect 25004 15524 25493 15552
rect 25004 15512 25010 15524
rect 25481 15521 25493 15524
rect 25527 15521 25539 15555
rect 27062 15552 27068 15564
rect 27023 15524 27068 15552
rect 25481 15515 25539 15521
rect 27062 15512 27068 15524
rect 27120 15512 27126 15564
rect 27246 15552 27252 15564
rect 27207 15524 27252 15552
rect 27246 15512 27252 15524
rect 27304 15512 27310 15564
rect 27430 15552 27436 15564
rect 27391 15524 27436 15552
rect 27430 15512 27436 15524
rect 27488 15512 27494 15564
rect 22557 15487 22615 15493
rect 22557 15453 22569 15487
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 25225 15487 25283 15493
rect 25225 15453 25237 15487
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 21361 15419 21419 15425
rect 21361 15385 21373 15419
rect 21407 15385 21419 15419
rect 22094 15416 22100 15428
rect 22055 15388 22100 15416
rect 21361 15379 21419 15385
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 20714 15348 20720 15360
rect 19996 15320 20720 15348
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22572 15348 22600 15447
rect 21968 15320 22600 15348
rect 25240 15348 25268 15447
rect 25406 15348 25412 15360
rect 25240 15320 25412 15348
rect 21968 15308 21974 15320
rect 25406 15308 25412 15320
rect 25464 15308 25470 15360
rect 26694 15308 26700 15360
rect 26752 15348 26758 15360
rect 27617 15351 27675 15357
rect 27617 15348 27629 15351
rect 26752 15320 27629 15348
rect 26752 15308 26758 15320
rect 27617 15317 27629 15320
rect 27663 15317 27675 15351
rect 27617 15311 27675 15317
rect 1104 15258 28428 15280
rect 1104 15206 5536 15258
rect 5588 15206 5600 15258
rect 5652 15206 5664 15258
rect 5716 15206 5728 15258
rect 5780 15206 14644 15258
rect 14696 15206 14708 15258
rect 14760 15206 14772 15258
rect 14824 15206 14836 15258
rect 14888 15206 23752 15258
rect 23804 15206 23816 15258
rect 23868 15206 23880 15258
rect 23932 15206 23944 15258
rect 23996 15206 28428 15258
rect 1104 15184 28428 15206
rect 4338 15144 4344 15156
rect 4299 15116 4344 15144
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 13078 15144 13084 15156
rect 7156 15116 13084 15144
rect 7156 15104 7162 15116
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 13354 15144 13360 15156
rect 13311 15116 13360 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 14458 15104 14464 15156
rect 14516 15144 14522 15156
rect 23198 15144 23204 15156
rect 14516 15116 23204 15144
rect 14516 15104 14522 15116
rect 23198 15104 23204 15116
rect 23256 15104 23262 15156
rect 23382 15144 23388 15156
rect 23343 15116 23388 15144
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24489 15147 24547 15153
rect 24489 15113 24501 15147
rect 24535 15144 24547 15147
rect 24854 15144 24860 15156
rect 24535 15116 24860 15144
rect 24535 15113 24547 15116
rect 24489 15107 24547 15113
rect 24854 15104 24860 15116
rect 24912 15104 24918 15156
rect 26881 15147 26939 15153
rect 26881 15113 26893 15147
rect 26927 15144 26939 15147
rect 27430 15144 27436 15156
rect 26927 15116 27436 15144
rect 26927 15113 26939 15116
rect 26881 15107 26939 15113
rect 27430 15104 27436 15116
rect 27488 15104 27494 15156
rect 9214 15036 9220 15088
rect 9272 15076 9278 15088
rect 9490 15076 9496 15088
rect 9272 15048 9496 15076
rect 9272 15036 9278 15048
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 9122 15008 9128 15020
rect 6972 14980 9128 15008
rect 6972 14968 6978 14980
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 2961 14943 3019 14949
rect 2961 14940 2973 14943
rect 2832 14912 2973 14940
rect 2832 14900 2838 14912
rect 2961 14909 2973 14912
rect 3007 14909 3019 14943
rect 2961 14903 3019 14909
rect 3228 14943 3286 14949
rect 3228 14909 3240 14943
rect 3274 14940 3286 14943
rect 4154 14940 4160 14952
rect 3274 14912 4160 14940
rect 3274 14909 3286 14912
rect 3228 14903 3286 14909
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 8294 14940 8300 14952
rect 8255 14912 8300 14940
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8754 14940 8760 14952
rect 8715 14912 8760 14940
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14909 9091 14943
rect 9306 14940 9312 14952
rect 9267 14912 9312 14940
rect 9033 14903 9091 14909
rect 8938 14872 8944 14884
rect 1596 14844 8944 14872
rect 1596 14813 1624 14844
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 9048 14872 9076 14903
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9416 14949 9444 15048
rect 9490 15036 9496 15048
rect 9548 15036 9554 15088
rect 9585 15079 9643 15085
rect 9585 15045 9597 15079
rect 9631 15045 9643 15079
rect 10686 15076 10692 15088
rect 10647 15048 10692 15076
rect 9585 15039 9643 15045
rect 9600 15008 9628 15039
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 15286 15076 15292 15088
rect 15247 15048 15292 15076
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 18506 15036 18512 15088
rect 18564 15076 18570 15088
rect 20254 15076 20260 15088
rect 18564 15048 19334 15076
rect 20215 15048 20260 15076
rect 18564 15036 18570 15048
rect 11330 15008 11336 15020
rect 9600 14980 11336 15008
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 11572 14980 12357 15008
rect 11572 14968 11578 14980
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 14090 14968 14096 15020
rect 14148 15008 14154 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14148 14980 14289 15008
rect 14148 14968 14154 14980
rect 14277 14977 14289 14980
rect 14323 15008 14335 15011
rect 14323 14980 15148 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 9732 14912 12173 14940
rect 9732 14900 9738 14912
rect 12161 14909 12173 14912
rect 12207 14940 12219 14943
rect 12207 14912 12572 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 10410 14872 10416 14884
rect 9048 14844 10416 14872
rect 10410 14832 10416 14844
rect 10468 14832 10474 14884
rect 10505 14875 10563 14881
rect 10505 14841 10517 14875
rect 10551 14872 10563 14875
rect 11422 14872 11428 14884
rect 10551 14844 11428 14872
rect 10551 14841 10563 14844
rect 10505 14835 10563 14841
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 12544 14872 12572 14912
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 12676 14912 13185 14940
rect 12676 14900 12682 14912
rect 13173 14909 13185 14912
rect 13219 14909 13231 14943
rect 14182 14940 14188 14952
rect 13173 14903 13231 14909
rect 14016 14912 14188 14940
rect 14016 14872 14044 14912
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14734 14940 14740 14952
rect 14695 14912 14740 14940
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 14918 14940 14924 14952
rect 14879 14912 14924 14940
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 15120 14949 15148 14980
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 17368 14980 17785 15008
rect 17368 14968 17374 14980
rect 17773 14977 17785 14980
rect 17819 15008 17831 15011
rect 17954 15008 17960 15020
rect 17819 14980 17960 15008
rect 17819 14977 17831 14980
rect 17773 14971 17831 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18782 15008 18788 15020
rect 18064 14980 18788 15008
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15286 14940 15292 14952
rect 15151 14912 15292 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 17497 14943 17555 14949
rect 17497 14909 17509 14943
rect 17543 14909 17555 14943
rect 17497 14903 17555 14909
rect 11808 14844 12368 14872
rect 12544 14844 14044 14872
rect 14093 14875 14151 14881
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 6917 14807 6975 14813
rect 6917 14773 6929 14807
rect 6963 14804 6975 14807
rect 7466 14804 7472 14816
rect 6963 14776 7472 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 7926 14764 7932 14816
rect 7984 14804 7990 14816
rect 11808 14804 11836 14844
rect 7984 14776 11836 14804
rect 12340 14804 12368 14844
rect 14093 14841 14105 14875
rect 14139 14872 14151 14875
rect 14826 14872 14832 14884
rect 14139 14844 14832 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15013 14875 15071 14881
rect 15013 14841 15025 14875
rect 15059 14872 15071 14875
rect 15746 14872 15752 14884
rect 15059 14844 15752 14872
rect 15059 14841 15071 14844
rect 15013 14835 15071 14841
rect 15746 14832 15752 14844
rect 15804 14832 15810 14884
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14872 15899 14875
rect 17512 14872 17540 14903
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 17865 14943 17923 14949
rect 17644 14912 17689 14940
rect 17644 14900 17650 14912
rect 17865 14909 17877 14943
rect 17911 14940 17923 14943
rect 18064 14940 18092 14980
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 17911 14912 18092 14940
rect 17911 14909 17923 14912
rect 17865 14903 17923 14909
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18380 14912 18521 14940
rect 18380 14900 18386 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 18874 14872 18880 14884
rect 15887 14844 17448 14872
rect 17512 14844 18880 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 14458 14804 14464 14816
rect 12340 14776 14464 14804
rect 7984 14764 7990 14776
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15933 14807 15991 14813
rect 15933 14804 15945 14807
rect 14792 14776 15945 14804
rect 14792 14764 14798 14776
rect 15933 14773 15945 14776
rect 15979 14773 15991 14807
rect 15933 14767 15991 14773
rect 16850 14764 16856 14816
rect 16908 14804 16914 14816
rect 17313 14807 17371 14813
rect 17313 14804 17325 14807
rect 16908 14776 17325 14804
rect 16908 14764 16914 14776
rect 17313 14773 17325 14776
rect 17359 14773 17371 14807
rect 17420 14804 17448 14844
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 19306 14872 19334 15048
rect 20254 15036 20260 15048
rect 20312 15036 20318 15088
rect 21634 15076 21640 15088
rect 21595 15048 21640 15076
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 23474 15076 23480 15088
rect 22152 15048 23480 15076
rect 22152 15036 22158 15048
rect 20916 14980 22416 15008
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 19705 14943 19763 14949
rect 19705 14940 19717 14943
rect 19576 14912 19717 14940
rect 19576 14900 19582 14912
rect 19705 14909 19717 14912
rect 19751 14909 19763 14943
rect 19886 14940 19892 14952
rect 19847 14912 19892 14940
rect 19705 14903 19763 14909
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 20070 14940 20076 14952
rect 20031 14912 20076 14940
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 19306 14844 19932 14872
rect 18322 14804 18328 14816
rect 17420 14776 18328 14804
rect 17313 14767 17371 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 18601 14807 18659 14813
rect 18601 14773 18613 14807
rect 18647 14804 18659 14807
rect 19702 14804 19708 14816
rect 18647 14776 19708 14804
rect 18647 14773 18659 14776
rect 18601 14767 18659 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 19904 14804 19932 14844
rect 19978 14832 19984 14884
rect 20036 14872 20042 14884
rect 20916 14872 20944 14980
rect 21082 14940 21088 14952
rect 21043 14912 21088 14940
rect 21082 14900 21088 14912
rect 21140 14900 21146 14952
rect 21266 14940 21272 14952
rect 21227 14912 21272 14940
rect 21266 14900 21272 14912
rect 21324 14900 21330 14952
rect 21453 14943 21511 14949
rect 21453 14909 21465 14943
rect 21499 14909 21511 14943
rect 21453 14903 21511 14909
rect 21358 14872 21364 14884
rect 20036 14844 20944 14872
rect 21319 14844 21364 14872
rect 20036 14832 20042 14844
rect 21358 14832 21364 14844
rect 21416 14832 21422 14884
rect 21468 14804 21496 14903
rect 22388 14872 22416 14980
rect 22833 14943 22891 14949
rect 22833 14909 22845 14943
rect 22879 14940 22891 14943
rect 22922 14940 22928 14952
rect 22879 14912 22928 14940
rect 22879 14909 22891 14912
rect 22833 14903 22891 14909
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 23032 14949 23060 15048
rect 23474 15036 23480 15048
rect 23532 15076 23538 15088
rect 23532 15048 24072 15076
rect 23532 15036 23538 15048
rect 23017 14943 23075 14949
rect 23017 14909 23029 14943
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14940 23259 14943
rect 23290 14940 23296 14952
rect 23247 14912 23296 14940
rect 23247 14909 23259 14912
rect 23201 14903 23259 14909
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23474 14900 23480 14952
rect 23532 14940 23538 14952
rect 23937 14943 23995 14949
rect 23937 14940 23949 14943
rect 23532 14912 23949 14940
rect 23532 14900 23538 14912
rect 23937 14909 23949 14912
rect 23983 14909 23995 14943
rect 23937 14903 23995 14909
rect 23109 14875 23167 14881
rect 23109 14872 23121 14875
rect 22388 14844 23121 14872
rect 23109 14841 23121 14844
rect 23155 14872 23167 14875
rect 23566 14872 23572 14884
rect 23155 14844 23572 14872
rect 23155 14841 23167 14844
rect 23109 14835 23167 14841
rect 23566 14832 23572 14844
rect 23624 14832 23630 14884
rect 24044 14872 24072 15048
rect 24210 14940 24216 14952
rect 24171 14912 24216 14940
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 24305 14943 24363 14949
rect 24305 14909 24317 14943
rect 24351 14940 24363 14943
rect 25222 14940 25228 14952
rect 24351 14912 25228 14940
rect 24351 14909 24363 14912
rect 24305 14903 24363 14909
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 25501 14943 25559 14949
rect 25501 14909 25513 14943
rect 25547 14909 25559 14943
rect 25501 14903 25559 14909
rect 25768 14943 25826 14949
rect 25768 14909 25780 14943
rect 25814 14940 25826 14943
rect 26694 14940 26700 14952
rect 25814 14912 26700 14940
rect 25814 14909 25826 14912
rect 25768 14903 25826 14909
rect 24121 14875 24179 14881
rect 24121 14872 24133 14875
rect 24044 14844 24133 14872
rect 24121 14841 24133 14844
rect 24167 14872 24179 14875
rect 24578 14872 24584 14884
rect 24167 14844 24584 14872
rect 24167 14841 24179 14844
rect 24121 14835 24179 14841
rect 24578 14832 24584 14844
rect 24636 14832 24642 14884
rect 25130 14832 25136 14884
rect 25188 14872 25194 14884
rect 25406 14872 25412 14884
rect 25188 14844 25412 14872
rect 25188 14832 25194 14844
rect 25406 14832 25412 14844
rect 25464 14872 25470 14884
rect 25516 14872 25544 14903
rect 26694 14900 26700 14912
rect 26752 14900 26758 14952
rect 26050 14872 26056 14884
rect 25464 14844 26056 14872
rect 25464 14832 25470 14844
rect 26050 14832 26056 14844
rect 26108 14832 26114 14884
rect 22462 14804 22468 14816
rect 19904 14776 22468 14804
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 1104 14714 28428 14736
rect 1104 14662 10090 14714
rect 10142 14662 10154 14714
rect 10206 14662 10218 14714
rect 10270 14662 10282 14714
rect 10334 14662 19198 14714
rect 19250 14662 19262 14714
rect 19314 14662 19326 14714
rect 19378 14662 19390 14714
rect 19442 14662 28428 14714
rect 1104 14640 28428 14662
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 8386 14600 8392 14612
rect 7156 14572 7236 14600
rect 7156 14560 7162 14572
rect 2406 14492 2412 14544
rect 2464 14532 2470 14544
rect 7208 14541 7236 14572
rect 7300 14572 8392 14600
rect 7300 14541 7328 14572
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 9398 14600 9404 14612
rect 8720 14572 9404 14600
rect 8720 14560 8726 14572
rect 9398 14560 9404 14572
rect 9456 14600 9462 14612
rect 9858 14600 9864 14612
rect 9456 14572 9864 14600
rect 9456 14560 9462 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 11054 14600 11060 14612
rect 10244 14572 11060 14600
rect 7193 14535 7251 14541
rect 2464 14504 7144 14532
rect 2464 14492 2470 14504
rect 1854 14464 1860 14476
rect 1815 14436 1860 14464
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 4338 14424 4344 14476
rect 4396 14464 4402 14476
rect 4709 14467 4767 14473
rect 4709 14464 4721 14467
rect 4396 14436 4721 14464
rect 4396 14424 4402 14436
rect 4709 14433 4721 14436
rect 4755 14433 4767 14467
rect 5902 14464 5908 14476
rect 5863 14436 5908 14464
rect 4709 14427 4767 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6012 14436 7021 14464
rect 1946 14356 1952 14408
rect 2004 14396 2010 14408
rect 6012 14396 6040 14436
rect 2004 14368 6040 14396
rect 6932 14396 6960 14436
rect 7009 14433 7021 14436
rect 7055 14433 7067 14467
rect 7116 14464 7144 14504
rect 7193 14501 7205 14535
rect 7239 14501 7251 14535
rect 7193 14495 7251 14501
rect 7285 14535 7343 14541
rect 7285 14501 7297 14535
rect 7331 14501 7343 14535
rect 9769 14535 9827 14541
rect 9769 14532 9781 14535
rect 7285 14495 7343 14501
rect 7392 14504 9781 14532
rect 7392 14473 7420 14504
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7116 14436 7389 14464
rect 7009 14427 7067 14433
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7650 14464 7656 14476
rect 7377 14427 7435 14433
rect 7484 14436 7656 14464
rect 7484 14396 7512 14436
rect 7650 14424 7656 14436
rect 7708 14464 7714 14476
rect 8404 14473 8432 14504
rect 9769 14501 9781 14504
rect 9815 14501 9827 14535
rect 9769 14495 9827 14501
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7708 14436 8033 14464
rect 7708 14424 7714 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14433 8263 14467
rect 8205 14427 8263 14433
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9674 14464 9680 14476
rect 9631 14436 9680 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 6932 14368 7512 14396
rect 2004 14356 2010 14368
rect 7834 14356 7840 14408
rect 7892 14396 7898 14408
rect 8220 14396 8248 14427
rect 7892 14368 8248 14396
rect 8312 14396 8340 14427
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10244 14473 10272 14572
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 22278 14600 22284 14612
rect 13372 14572 22284 14600
rect 10505 14535 10563 14541
rect 10505 14501 10517 14535
rect 10551 14532 10563 14535
rect 10870 14532 10876 14544
rect 10551 14504 10876 14532
rect 10551 14501 10563 14504
rect 10505 14495 10563 14501
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14433 10287 14467
rect 10410 14464 10416 14476
rect 10371 14436 10416 14464
rect 10229 14427 10287 14433
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 10962 14464 10968 14476
rect 10643 14436 10968 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 11497 14467 11555 14473
rect 11497 14464 11509 14467
rect 11204 14436 11509 14464
rect 11204 14424 11210 14436
rect 11497 14433 11509 14436
rect 11543 14433 11555 14467
rect 11497 14427 11555 14433
rect 8312 14368 8432 14396
rect 7892 14356 7898 14368
rect 2038 14328 2044 14340
rect 1999 14300 2044 14328
rect 2038 14288 2044 14300
rect 2096 14288 2102 14340
rect 5169 14331 5227 14337
rect 5169 14297 5181 14331
rect 5215 14328 5227 14331
rect 6730 14328 6736 14340
rect 5215 14300 6736 14328
rect 5215 14297 5227 14300
rect 5169 14291 5227 14297
rect 6730 14288 6736 14300
rect 6788 14288 6794 14340
rect 4985 14263 5043 14269
rect 4985 14229 4997 14263
rect 5031 14260 5043 14263
rect 5074 14260 5080 14272
rect 5031 14232 5080 14260
rect 5031 14229 5043 14232
rect 4985 14223 5043 14229
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5408 14232 6009 14260
rect 5408 14220 5414 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 5997 14223 6055 14229
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7650 14260 7656 14272
rect 7607 14232 7656 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8404 14260 8432 14368
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 10778 14396 10784 14408
rect 9180 14368 10784 14396
rect 9180 14356 9186 14368
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11238 14396 11244 14408
rect 11199 14368 11244 14396
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 13372 14328 13400 14572
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 22373 14603 22431 14609
rect 22373 14569 22385 14603
rect 22419 14600 22431 14603
rect 22462 14600 22468 14612
rect 22419 14572 22468 14600
rect 22419 14569 22431 14572
rect 22373 14563 22431 14569
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 25869 14603 25927 14609
rect 25869 14569 25881 14603
rect 25915 14569 25927 14603
rect 25869 14563 25927 14569
rect 15010 14532 15016 14544
rect 14923 14504 15016 14532
rect 15010 14492 15016 14504
rect 15068 14532 15074 14544
rect 15930 14532 15936 14544
rect 15068 14504 15936 14532
rect 15068 14492 15074 14504
rect 15930 14492 15936 14504
rect 15988 14492 15994 14544
rect 16298 14492 16304 14544
rect 16356 14532 16362 14544
rect 16393 14535 16451 14541
rect 16393 14532 16405 14535
rect 16356 14504 16405 14532
rect 16356 14492 16362 14504
rect 16393 14501 16405 14504
rect 16439 14501 16451 14535
rect 16393 14495 16451 14501
rect 16758 14492 16764 14544
rect 16816 14532 16822 14544
rect 16816 14504 17172 14532
rect 16816 14492 16822 14504
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13630 14464 13636 14476
rect 13504 14436 13636 14464
rect 13504 14424 13510 14436
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 14734 14464 14740 14476
rect 14695 14436 14740 14464
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 14918 14464 14924 14476
rect 14835 14436 14924 14464
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14835 14396 14863 14436
rect 14918 14424 14924 14436
rect 14976 14424 14982 14476
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14464 15163 14467
rect 15286 14464 15292 14476
rect 15151 14436 15292 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 16114 14464 16120 14476
rect 15712 14436 16120 14464
rect 15712 14424 15718 14436
rect 16114 14424 16120 14436
rect 16172 14464 16178 14476
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 16172 14436 16221 14464
rect 16172 14424 16178 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 16850 14464 16856 14476
rect 16811 14436 16856 14464
rect 16209 14427 16267 14433
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 17144 14473 17172 14504
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 19610 14532 19616 14544
rect 18380 14504 19616 14532
rect 18380 14492 18386 14504
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 21260 14535 21318 14541
rect 21260 14501 21272 14535
rect 21306 14532 21318 14535
rect 21634 14532 21640 14544
rect 21306 14504 21640 14532
rect 21306 14501 21318 14504
rect 21260 14495 21318 14501
rect 21634 14492 21640 14504
rect 21692 14492 21698 14544
rect 25590 14532 25596 14544
rect 25551 14504 25596 14532
rect 25590 14492 25596 14504
rect 25648 14492 25654 14544
rect 25884 14532 25912 14563
rect 26574 14535 26632 14541
rect 26574 14532 26586 14535
rect 25884 14504 26586 14532
rect 26574 14501 26586 14504
rect 26620 14501 26632 14535
rect 26574 14495 26632 14501
rect 17037 14467 17095 14473
rect 17037 14433 17049 14467
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 17132 14467 17190 14473
rect 17132 14433 17144 14467
rect 17178 14433 17190 14467
rect 17132 14427 17190 14433
rect 14516 14368 14863 14396
rect 17052 14396 17080 14427
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 17402 14464 17408 14476
rect 17276 14436 17321 14464
rect 17363 14436 17408 14464
rect 17276 14424 17282 14436
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18046 14464 18052 14476
rect 17512 14436 18052 14464
rect 17512 14396 17540 14436
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14464 18199 14467
rect 18506 14464 18512 14476
rect 18187 14436 18512 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 20073 14467 20131 14473
rect 20073 14433 20085 14467
rect 20119 14464 20131 14467
rect 20622 14464 20628 14476
rect 20119 14436 20628 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 20993 14467 21051 14473
rect 20993 14464 21005 14467
rect 20772 14436 21005 14464
rect 20772 14424 20778 14436
rect 20993 14433 21005 14436
rect 21039 14464 21051 14467
rect 21818 14464 21824 14476
rect 21039 14436 21824 14464
rect 21039 14433 21051 14436
rect 20993 14427 21051 14433
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 23198 14424 23204 14476
rect 23256 14464 23262 14476
rect 25317 14467 25375 14473
rect 25317 14464 25329 14467
rect 23256 14436 25329 14464
rect 23256 14424 23262 14436
rect 25317 14433 25329 14436
rect 25363 14433 25375 14467
rect 25498 14464 25504 14476
rect 25459 14436 25504 14464
rect 25317 14427 25375 14433
rect 25498 14424 25504 14436
rect 25556 14424 25562 14476
rect 25685 14467 25743 14473
rect 25685 14433 25697 14467
rect 25731 14464 25743 14467
rect 27430 14464 27436 14476
rect 25731 14436 27436 14464
rect 25731 14433 25743 14436
rect 25685 14427 25743 14433
rect 27430 14424 27436 14436
rect 27488 14464 27494 14476
rect 27488 14436 27752 14464
rect 27488 14424 27494 14436
rect 17052 14368 17540 14396
rect 17589 14399 17647 14405
rect 14516 14356 14522 14368
rect 17589 14365 17601 14399
rect 17635 14396 17647 14399
rect 18874 14396 18880 14408
rect 17635 14368 18880 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 18966 14356 18972 14408
rect 19024 14396 19030 14408
rect 20806 14396 20812 14408
rect 19024 14368 20812 14396
rect 19024 14356 19030 14368
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 26329 14399 26387 14405
rect 26329 14365 26341 14399
rect 26375 14365 26387 14399
rect 26329 14359 26387 14365
rect 8628 14300 11284 14328
rect 8628 14288 8634 14300
rect 8662 14260 8668 14272
rect 8404 14232 8668 14260
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 9950 14260 9956 14272
rect 8996 14232 9956 14260
rect 8996 14220 9002 14232
rect 9950 14220 9956 14232
rect 10008 14260 10014 14272
rect 10410 14260 10416 14272
rect 10008 14232 10416 14260
rect 10008 14220 10014 14232
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 10778 14260 10784 14272
rect 10739 14232 10784 14260
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11256 14260 11284 14300
rect 12176 14300 13400 14328
rect 12176 14260 12204 14300
rect 13446 14288 13452 14340
rect 13504 14328 13510 14340
rect 20257 14331 20315 14337
rect 13504 14300 19334 14328
rect 13504 14288 13510 14300
rect 11256 14232 12204 14260
rect 12621 14263 12679 14269
rect 12621 14229 12633 14263
rect 12667 14260 12679 14263
rect 12986 14260 12992 14272
rect 12667 14232 12992 14260
rect 12667 14229 12679 14232
rect 12621 14223 12679 14229
rect 12986 14220 12992 14232
rect 13044 14220 13050 14272
rect 13722 14260 13728 14272
rect 13683 14232 13728 14260
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 15252 14232 15301 14260
rect 15252 14220 15258 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 15289 14223 15347 14229
rect 17494 14220 17500 14272
rect 17552 14260 17558 14272
rect 18046 14260 18052 14272
rect 17552 14232 18052 14260
rect 17552 14220 17558 14232
rect 18046 14220 18052 14232
rect 18104 14260 18110 14272
rect 18233 14263 18291 14269
rect 18233 14260 18245 14263
rect 18104 14232 18245 14260
rect 18104 14220 18110 14232
rect 18233 14229 18245 14232
rect 18279 14229 18291 14263
rect 19306 14260 19334 14300
rect 20257 14297 20269 14331
rect 20303 14328 20315 14331
rect 20530 14328 20536 14340
rect 20303 14300 20536 14328
rect 20303 14297 20315 14300
rect 20257 14291 20315 14297
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 23106 14288 23112 14340
rect 23164 14328 23170 14340
rect 23164 14300 25912 14328
rect 23164 14288 23170 14300
rect 25774 14260 25780 14272
rect 19306 14232 25780 14260
rect 18233 14223 18291 14229
rect 25774 14220 25780 14232
rect 25832 14220 25838 14272
rect 25884 14260 25912 14300
rect 26050 14288 26056 14340
rect 26108 14328 26114 14340
rect 26344 14328 26372 14359
rect 27724 14337 27752 14436
rect 26108 14300 26372 14328
rect 27709 14331 27767 14337
rect 26108 14288 26114 14300
rect 27709 14297 27721 14331
rect 27755 14297 27767 14331
rect 27709 14291 27767 14297
rect 27062 14260 27068 14272
rect 25884 14232 27068 14260
rect 27062 14220 27068 14232
rect 27120 14220 27126 14272
rect 1104 14170 28428 14192
rect 1104 14118 5536 14170
rect 5588 14118 5600 14170
rect 5652 14118 5664 14170
rect 5716 14118 5728 14170
rect 5780 14118 14644 14170
rect 14696 14118 14708 14170
rect 14760 14118 14772 14170
rect 14824 14118 14836 14170
rect 14888 14118 23752 14170
rect 23804 14118 23816 14170
rect 23868 14118 23880 14170
rect 23932 14118 23944 14170
rect 23996 14118 28428 14170
rect 1104 14096 28428 14118
rect 7098 14056 7104 14068
rect 5552 14028 7104 14056
rect 5552 14000 5580 14028
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8941 14059 8999 14065
rect 8941 14056 8953 14059
rect 8536 14028 8953 14056
rect 8536 14016 8542 14028
rect 8941 14025 8953 14028
rect 8987 14025 8999 14059
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 8941 14019 8999 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 23106 14056 23112 14068
rect 11388 14028 23112 14056
rect 11388 14016 11394 14028
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23198 14016 23204 14068
rect 23256 14056 23262 14068
rect 24946 14056 24952 14068
rect 23256 14028 23520 14056
rect 24907 14028 24952 14056
rect 23256 14016 23262 14028
rect 3421 13991 3479 13997
rect 3421 13957 3433 13991
rect 3467 13988 3479 13991
rect 4338 13988 4344 14000
rect 3467 13960 4344 13988
rect 3467 13957 3479 13960
rect 3421 13951 3479 13957
rect 4338 13948 4344 13960
rect 4396 13988 4402 14000
rect 5350 13988 5356 14000
rect 4396 13960 5356 13988
rect 4396 13948 4402 13960
rect 5350 13948 5356 13960
rect 5408 13948 5414 14000
rect 5534 13948 5540 14000
rect 5592 13948 5598 14000
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 11054 13988 11060 14000
rect 6696 13960 7604 13988
rect 6696 13948 6702 13960
rect 3234 13920 3240 13932
rect 2148 13892 3240 13920
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2148 13861 2176 13892
rect 3234 13880 3240 13892
rect 3292 13920 3298 13932
rect 4982 13920 4988 13932
rect 3292 13892 3740 13920
rect 3292 13880 3298 13892
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13821 2191 13855
rect 2133 13815 2191 13821
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2406 13852 2412 13864
rect 2363 13824 2412 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 3712 13861 3740 13892
rect 3896 13892 4988 13920
rect 3896 13861 3924 13892
rect 4982 13880 4988 13892
rect 5040 13920 5046 13932
rect 5040 13892 5764 13920
rect 5040 13880 5046 13892
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 3467 13824 3525 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 3513 13821 3525 13824
rect 3559 13821 3571 13855
rect 3513 13815 3571 13821
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 3881 13855 3939 13861
rect 3881 13821 3893 13855
rect 3927 13821 3939 13855
rect 5350 13852 5356 13864
rect 5311 13824 5356 13852
rect 3881 13815 3939 13821
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5534 13852 5540 13864
rect 5495 13824 5540 13852
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5736 13861 5764 13892
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 7576 13929 7604 13960
rect 10612 13960 11060 13988
rect 7561 13923 7619 13929
rect 5960 13892 7512 13920
rect 5960 13880 5966 13892
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 5767 13824 7113 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 2222 13784 2228 13796
rect 2183 13756 2228 13784
rect 2222 13744 2228 13756
rect 2280 13744 2286 13796
rect 3789 13787 3847 13793
rect 3789 13753 3801 13787
rect 3835 13784 3847 13787
rect 4246 13784 4252 13796
rect 3835 13756 4252 13784
rect 3835 13753 3847 13756
rect 3789 13747 3847 13753
rect 4246 13744 4252 13756
rect 4304 13744 4310 13796
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13784 5687 13787
rect 6822 13784 6828 13796
rect 5675 13756 6828 13784
rect 5675 13753 5687 13756
rect 5629 13747 5687 13753
rect 6822 13744 6828 13756
rect 6880 13744 6886 13796
rect 6914 13744 6920 13796
rect 6972 13784 6978 13796
rect 7484 13784 7512 13892
rect 7561 13889 7573 13923
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 7817 13855 7875 13861
rect 7817 13852 7829 13855
rect 7708 13824 7829 13852
rect 7708 13812 7714 13824
rect 7817 13821 7829 13824
rect 7863 13821 7875 13855
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 7817 13815 7875 13821
rect 7944 13824 9965 13852
rect 7944 13784 7972 13824
rect 9953 13821 9965 13824
rect 9999 13852 10011 13855
rect 10318 13852 10324 13864
rect 9999 13824 10324 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10612 13861 10640 13960
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 13446 13988 13452 14000
rect 13407 13960 13452 13988
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 14182 13948 14188 14000
rect 14240 13988 14246 14000
rect 14277 13991 14335 13997
rect 14277 13988 14289 13991
rect 14240 13960 14289 13988
rect 14240 13948 14246 13960
rect 14277 13957 14289 13960
rect 14323 13957 14335 13991
rect 14277 13951 14335 13957
rect 20533 13991 20591 13997
rect 20533 13957 20545 13991
rect 20579 13988 20591 13991
rect 20579 13960 23428 13988
rect 20579 13957 20591 13960
rect 20533 13951 20591 13957
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 16022 13920 16028 13932
rect 13136 13892 14863 13920
rect 15983 13892 16028 13920
rect 13136 13880 13142 13892
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13821 10655 13855
rect 10778 13852 10784 13864
rect 10739 13824 10784 13852
rect 10597 13815 10655 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 10962 13852 10968 13864
rect 10875 13824 10968 13852
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 11330 13812 11336 13864
rect 11388 13852 11394 13864
rect 12066 13852 12072 13864
rect 11388 13824 12072 13852
rect 11388 13812 11394 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12325 13855 12383 13861
rect 12325 13852 12337 13855
rect 12216 13824 12337 13852
rect 12216 13812 12222 13824
rect 12325 13821 12337 13824
rect 12371 13821 12383 13855
rect 12325 13815 12383 13821
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14366 13852 14372 13864
rect 13964 13824 14372 13852
rect 13964 13812 13970 13824
rect 14366 13812 14372 13824
rect 14424 13852 14430 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14424 13824 14749 13852
rect 14424 13812 14430 13824
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 14835 13852 14863 13892
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 19702 13880 19708 13932
rect 19760 13920 19766 13932
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19760 13892 19993 13920
rect 19760 13880 19766 13892
rect 19981 13889 19993 13892
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 20128 13892 20760 13920
rect 20128 13880 20134 13892
rect 15102 13852 15108 13864
rect 15160 13861 15166 13864
rect 15160 13855 15187 13861
rect 14835 13824 15108 13852
rect 14737 13815 14795 13821
rect 15102 13812 15108 13824
rect 15175 13821 15187 13855
rect 15160 13815 15187 13821
rect 15160 13812 15166 13815
rect 17034 13812 17040 13864
rect 17092 13852 17098 13864
rect 17865 13855 17923 13861
rect 17865 13852 17877 13855
rect 17092 13824 17877 13852
rect 17092 13812 17098 13824
rect 17865 13821 17877 13824
rect 17911 13821 17923 13855
rect 17865 13815 17923 13821
rect 18874 13812 18880 13864
rect 18932 13852 18938 13864
rect 19797 13855 19855 13861
rect 19797 13852 19809 13855
rect 18932 13824 19809 13852
rect 18932 13812 18938 13824
rect 19797 13821 19809 13824
rect 19843 13821 19855 13855
rect 20254 13852 20260 13864
rect 20215 13824 20260 13852
rect 19797 13815 19855 13821
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 20622 13852 20628 13864
rect 20583 13824 20628 13852
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 20732 13861 20760 13892
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 20898 13812 20904 13864
rect 20956 13852 20962 13864
rect 23400 13861 23428 13960
rect 23492 13920 23520 14028
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 25682 14016 25688 14068
rect 25740 14056 25746 14068
rect 26050 14056 26056 14068
rect 25740 14028 26056 14056
rect 25740 14016 25746 14028
rect 26050 14016 26056 14028
rect 26108 14016 26114 14068
rect 23937 13991 23995 13997
rect 23937 13957 23949 13991
rect 23983 13988 23995 13991
rect 25406 13988 25412 14000
rect 23983 13960 25412 13988
rect 23983 13957 23995 13960
rect 23937 13951 23995 13957
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 26142 13988 26148 14000
rect 26103 13960 26148 13988
rect 26142 13948 26148 13960
rect 26200 13948 26206 14000
rect 26510 13920 26516 13932
rect 23492 13892 24440 13920
rect 21361 13855 21419 13861
rect 21361 13852 21373 13855
rect 20956 13824 21373 13852
rect 20956 13812 20962 13824
rect 21361 13821 21373 13824
rect 21407 13821 21419 13855
rect 21361 13815 21419 13821
rect 23385 13855 23443 13861
rect 23385 13821 23397 13855
rect 23431 13821 23443 13855
rect 23569 13855 23627 13861
rect 23569 13852 23581 13855
rect 23385 13815 23443 13821
rect 23492 13824 23581 13852
rect 6972 13756 7017 13784
rect 7484 13756 7972 13784
rect 10137 13787 10195 13793
rect 6972 13744 6978 13756
rect 10137 13753 10149 13787
rect 10183 13784 10195 13787
rect 10686 13784 10692 13796
rect 10183 13756 10692 13784
rect 10183 13753 10195 13756
rect 10137 13747 10195 13753
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 10873 13787 10931 13793
rect 10873 13753 10885 13787
rect 10919 13753 10931 13787
rect 10980 13784 11008 13812
rect 11514 13784 11520 13796
rect 10980 13756 11520 13784
rect 10873 13747 10931 13753
rect 2498 13716 2504 13728
rect 2459 13688 2504 13716
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 4062 13716 4068 13728
rect 4023 13688 4068 13716
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 5902 13716 5908 13728
rect 5863 13688 5908 13716
rect 5902 13676 5908 13688
rect 5960 13676 5966 13728
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 10888 13716 10916 13747
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 14093 13787 14151 13793
rect 14093 13753 14105 13787
rect 14139 13784 14151 13787
rect 14274 13784 14280 13796
rect 14139 13756 14280 13784
rect 14139 13753 14151 13756
rect 14093 13747 14151 13753
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 14516 13756 14933 13784
rect 14516 13744 14522 13756
rect 14921 13753 14933 13756
rect 14967 13753 14979 13787
rect 14921 13747 14979 13753
rect 15013 13787 15071 13793
rect 15013 13753 15025 13787
rect 15059 13784 15071 13787
rect 15562 13784 15568 13796
rect 15059 13756 15568 13784
rect 15059 13753 15071 13756
rect 15013 13747 15071 13753
rect 12986 13716 12992 13728
rect 6052 13688 12992 13716
rect 6052 13676 6058 13688
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 14936 13716 14964 13747
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 15841 13787 15899 13793
rect 15841 13753 15853 13787
rect 15887 13784 15899 13787
rect 16482 13784 16488 13796
rect 15887 13756 16488 13784
rect 15887 13753 15899 13756
rect 15841 13747 15899 13753
rect 16482 13744 16488 13756
rect 16540 13744 16546 13796
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 18110 13787 18168 13793
rect 18110 13784 18122 13787
rect 18012 13756 18122 13784
rect 18012 13744 18018 13756
rect 18110 13753 18122 13756
rect 18156 13753 18168 13787
rect 18110 13747 18168 13753
rect 18322 13744 18328 13796
rect 18380 13784 18386 13796
rect 20990 13784 20996 13796
rect 18380 13756 20996 13784
rect 18380 13744 18386 13756
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 23492 13784 23520 13824
rect 23569 13821 23581 13824
rect 23615 13821 23627 13855
rect 23569 13815 23627 13821
rect 23753 13855 23811 13861
rect 23753 13821 23765 13855
rect 23799 13852 23811 13855
rect 24302 13852 24308 13864
rect 23799 13824 24308 13852
rect 23799 13821 23811 13824
rect 23753 13815 23811 13821
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 24412 13861 24440 13892
rect 24780 13892 26516 13920
rect 24397 13855 24455 13861
rect 24397 13821 24409 13855
rect 24443 13821 24455 13855
rect 24578 13852 24584 13864
rect 24539 13824 24584 13852
rect 24397 13815 24455 13821
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 24780 13861 24808 13892
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 24765 13855 24823 13861
rect 24765 13821 24777 13855
rect 24811 13821 24823 13855
rect 24765 13815 24823 13821
rect 25774 13812 25780 13864
rect 25832 13852 25838 13864
rect 25961 13855 26019 13861
rect 25961 13852 25973 13855
rect 25832 13824 25973 13852
rect 25832 13812 25838 13824
rect 25961 13821 25973 13824
rect 26007 13852 26019 13855
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 26007 13824 26617 13852
rect 26007 13821 26019 13824
rect 25961 13815 26019 13821
rect 26605 13821 26617 13824
rect 26651 13821 26663 13855
rect 26605 13815 26663 13821
rect 23658 13784 23664 13796
rect 23400 13756 23520 13784
rect 23619 13756 23664 13784
rect 23400 13728 23428 13756
rect 23658 13744 23664 13756
rect 23716 13744 23722 13796
rect 24673 13787 24731 13793
rect 24673 13753 24685 13787
rect 24719 13753 24731 13787
rect 24673 13747 24731 13753
rect 15102 13716 15108 13728
rect 14936 13688 15108 13716
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15286 13716 15292 13728
rect 15247 13688 15292 13716
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 19058 13676 19064 13728
rect 19116 13716 19122 13728
rect 19245 13719 19303 13725
rect 19245 13716 19257 13719
rect 19116 13688 19257 13716
rect 19116 13676 19122 13688
rect 19245 13685 19257 13688
rect 19291 13685 19303 13719
rect 19245 13679 19303 13685
rect 20898 13676 20904 13728
rect 20956 13716 20962 13728
rect 21453 13719 21511 13725
rect 21453 13716 21465 13719
rect 20956 13688 21465 13716
rect 20956 13676 20962 13688
rect 21453 13685 21465 13688
rect 21499 13685 21511 13719
rect 21453 13679 21511 13685
rect 23382 13676 23388 13728
rect 23440 13676 23446 13728
rect 23676 13716 23704 13744
rect 24688 13716 24716 13747
rect 23676 13688 24716 13716
rect 1104 13626 28428 13648
rect 1104 13574 10090 13626
rect 10142 13574 10154 13626
rect 10206 13574 10218 13626
rect 10270 13574 10282 13626
rect 10334 13574 19198 13626
rect 19250 13574 19262 13626
rect 19314 13574 19326 13626
rect 19378 13574 19390 13626
rect 19442 13574 28428 13626
rect 1104 13552 28428 13574
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2280 13484 2881 13512
rect 2280 13472 2286 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 1756 13447 1814 13453
rect 1756 13413 1768 13447
rect 1802 13444 1814 13447
rect 2498 13444 2504 13456
rect 1802 13416 2504 13444
rect 1802 13413 1814 13416
rect 1756 13407 1814 13413
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 2884 13376 2912 13475
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 5074 13512 5080 13524
rect 4212 13484 5080 13512
rect 4212 13472 4218 13484
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 6822 13512 6828 13524
rect 6595 13484 6828 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13512 7343 13515
rect 8294 13512 8300 13524
rect 7331 13484 8300 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 9306 13512 9312 13524
rect 8435 13484 9312 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 10594 13512 10600 13524
rect 9723 13484 10600 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 10781 13515 10839 13521
rect 10781 13481 10793 13515
rect 10827 13481 10839 13515
rect 12618 13512 12624 13524
rect 10781 13475 10839 13481
rect 12406 13484 12624 13512
rect 5436 13447 5494 13453
rect 5436 13413 5448 13447
rect 5482 13444 5494 13447
rect 5902 13444 5908 13456
rect 5482 13416 5908 13444
rect 5482 13413 5494 13416
rect 5436 13407 5494 13413
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 9582 13444 9588 13456
rect 6012 13416 8432 13444
rect 9543 13416 9588 13444
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 2884 13348 4261 13376
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 5074 13336 5080 13388
rect 5132 13376 5138 13388
rect 6012 13376 6040 13416
rect 7466 13376 7472 13388
rect 5132 13348 6040 13376
rect 7427 13348 7472 13376
rect 5132 13336 5138 13348
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 7650 13376 7656 13388
rect 7607 13348 7656 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 7837 13339 7895 13345
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13277 1547 13311
rect 1489 13271 1547 13277
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 1504 13172 1532 13271
rect 5184 13240 5212 13271
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7852 13308 7880 13339
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8404 13376 8432 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 10505 13447 10563 13453
rect 10505 13413 10517 13447
rect 10551 13444 10563 13447
rect 10796 13444 10824 13475
rect 11486 13447 11544 13453
rect 11486 13444 11498 13447
rect 10551 13416 10732 13444
rect 10796 13416 11498 13444
rect 10551 13413 10563 13416
rect 10505 13407 10563 13413
rect 9766 13376 9772 13388
rect 8404 13348 9772 13376
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10410 13376 10416 13388
rect 10371 13348 10416 13376
rect 10229 13339 10287 13345
rect 6972 13280 7880 13308
rect 10244 13308 10272 13339
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 10594 13376 10600 13388
rect 10555 13348 10600 13376
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 10704 13376 10732 13416
rect 11486 13413 11498 13416
rect 11532 13413 11544 13447
rect 11486 13407 11544 13413
rect 12406 13376 12434 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 15160 13484 15323 13512
rect 15160 13472 15166 13484
rect 15004 13447 15062 13453
rect 15004 13413 15016 13447
rect 15050 13444 15062 13447
rect 15194 13444 15200 13456
rect 15050 13416 15200 13444
rect 15050 13413 15062 13416
rect 15004 13407 15062 13413
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 15295 13444 15323 13484
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15988 13484 16129 13512
rect 15988 13472 15994 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 17681 13515 17739 13521
rect 16117 13475 16175 13481
rect 16224 13484 17356 13512
rect 16224 13444 16252 13484
rect 15295 13416 16252 13444
rect 16298 13404 16304 13456
rect 16356 13444 16362 13456
rect 17328 13453 17356 13484
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 17954 13512 17960 13524
rect 17727 13484 17960 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 18966 13472 18972 13524
rect 19024 13512 19030 13524
rect 19024 13484 23796 13512
rect 19024 13472 19030 13484
rect 17313 13447 17371 13453
rect 16356 13416 17172 13444
rect 16356 13404 16362 13416
rect 10704 13348 12434 13376
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 17034 13376 17040 13388
rect 14783 13348 17040 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 17144 13385 17172 13416
rect 17313 13413 17325 13447
rect 17359 13413 17371 13447
rect 17313 13407 17371 13413
rect 17405 13447 17463 13453
rect 17405 13413 17417 13447
rect 17451 13444 17463 13447
rect 19058 13444 19064 13456
rect 17451 13416 19064 13444
rect 17451 13413 17463 13416
rect 17405 13407 17463 13413
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 21082 13444 21088 13456
rect 21043 13416 21088 13444
rect 21082 13404 21088 13416
rect 21140 13404 21146 13456
rect 17129 13379 17187 13385
rect 17129 13345 17141 13379
rect 17175 13345 17187 13379
rect 17129 13339 17187 13345
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 18230 13376 18236 13388
rect 18191 13348 18236 13376
rect 17497 13339 17555 13345
rect 10686 13308 10692 13320
rect 10244 13280 10692 13308
rect 6972 13268 6978 13280
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 11238 13308 11244 13320
rect 11199 13280 11244 13308
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17512 13308 17540 13339
rect 18230 13336 18236 13348
rect 18288 13336 18294 13388
rect 18874 13376 18880 13388
rect 18835 13348 18880 13376
rect 18874 13336 18880 13348
rect 18932 13336 18938 13388
rect 20073 13379 20131 13385
rect 20073 13345 20085 13379
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 20993 13379 21051 13385
rect 20993 13345 21005 13379
rect 21039 13376 21051 13379
rect 21453 13379 21511 13385
rect 21039 13348 21128 13376
rect 21039 13345 21051 13348
rect 20993 13339 21051 13345
rect 17368 13280 17540 13308
rect 17368 13268 17374 13280
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 20088 13308 20116 13339
rect 21100 13320 21128 13348
rect 21453 13345 21465 13379
rect 21499 13345 21511 13379
rect 21560 13376 21588 13484
rect 22557 13447 22615 13453
rect 22557 13444 22569 13447
rect 22020 13416 22569 13444
rect 22020 13385 22048 13416
rect 22557 13413 22569 13416
rect 22603 13413 22615 13447
rect 22557 13407 22615 13413
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21560 13348 21833 13376
rect 21453 13339 21511 13345
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 22005 13379 22063 13385
rect 22005 13345 22017 13379
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 18656 13280 20116 13308
rect 18656 13268 18662 13280
rect 21082 13268 21088 13320
rect 21140 13268 21146 13320
rect 4264 13212 5212 13240
rect 2774 13172 2780 13184
rect 1504 13144 2780 13172
rect 2774 13132 2780 13144
rect 2832 13172 2838 13184
rect 4264 13172 4292 13212
rect 2832 13144 4292 13172
rect 4341 13175 4399 13181
rect 2832 13132 2838 13144
rect 4341 13141 4353 13175
rect 4387 13172 4399 13175
rect 5074 13172 5080 13184
rect 4387 13144 5080 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5184 13172 5212 13212
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 7466 13240 7472 13252
rect 7340 13212 7472 13240
rect 7340 13200 7346 13212
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 7745 13243 7803 13249
rect 7745 13209 7757 13243
rect 7791 13240 7803 13243
rect 9030 13240 9036 13252
rect 7791 13212 9036 13240
rect 7791 13209 7803 13212
rect 7745 13203 7803 13209
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10778 13240 10784 13252
rect 10468 13212 10784 13240
rect 10468 13200 10474 13212
rect 10778 13200 10784 13212
rect 10836 13240 10842 13252
rect 10836 13212 11100 13240
rect 10836 13200 10842 13212
rect 6638 13172 6644 13184
rect 5184 13144 6644 13172
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 10962 13172 10968 13184
rect 7708 13144 10968 13172
rect 7708 13132 7714 13144
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11072 13172 11100 13212
rect 18046 13200 18052 13252
rect 18104 13240 18110 13252
rect 18966 13240 18972 13252
rect 18104 13212 18552 13240
rect 18927 13212 18972 13240
rect 18104 13200 18110 13212
rect 11606 13172 11612 13184
rect 11072 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 15930 13172 15936 13184
rect 13780 13144 15936 13172
rect 13780 13132 13786 13144
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 16666 13132 16672 13184
rect 16724 13172 16730 13184
rect 17678 13172 17684 13184
rect 16724 13144 17684 13172
rect 16724 13132 16730 13144
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 18325 13175 18383 13181
rect 18325 13141 18337 13175
rect 18371 13172 18383 13175
rect 18414 13172 18420 13184
rect 18371 13144 18420 13172
rect 18371 13141 18383 13144
rect 18325 13135 18383 13141
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 18524 13172 18552 13212
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 20257 13243 20315 13249
rect 20257 13209 20269 13243
rect 20303 13240 20315 13243
rect 20806 13240 20812 13252
rect 20303 13212 20812 13240
rect 20303 13209 20315 13212
rect 20257 13203 20315 13209
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 21468 13172 21496 13339
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 22465 13379 22523 13385
rect 22465 13376 22477 13379
rect 22152 13348 22477 13376
rect 22152 13336 22158 13348
rect 22465 13345 22477 13348
rect 22511 13345 22523 13379
rect 22465 13339 22523 13345
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13376 23259 13379
rect 23290 13376 23296 13388
rect 23247 13348 23296 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 23661 13379 23719 13385
rect 23661 13345 23673 13379
rect 23707 13345 23719 13379
rect 23768 13376 23796 13484
rect 24302 13472 24308 13524
rect 24360 13512 24366 13524
rect 25222 13512 25228 13524
rect 24360 13484 25228 13512
rect 24360 13472 24366 13484
rect 25222 13472 25228 13484
rect 25280 13512 25286 13524
rect 26605 13515 26663 13521
rect 26605 13512 26617 13515
rect 25280 13484 26617 13512
rect 25280 13472 25286 13484
rect 26605 13481 26617 13484
rect 26651 13481 26663 13515
rect 26605 13475 26663 13481
rect 25406 13404 25412 13456
rect 25464 13453 25470 13456
rect 25464 13447 25528 13453
rect 25464 13413 25482 13447
rect 25516 13413 25528 13447
rect 25464 13407 25528 13413
rect 25464 13404 25470 13407
rect 24029 13379 24087 13385
rect 24029 13376 24041 13379
rect 23768 13348 24041 13376
rect 23661 13339 23719 13345
rect 24029 13345 24041 13348
rect 24075 13376 24087 13379
rect 24118 13376 24124 13388
rect 24075 13348 24124 13376
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13277 21603 13311
rect 22554 13308 22560 13320
rect 21545 13271 21603 13277
rect 21836 13280 22560 13308
rect 21560 13240 21588 13271
rect 21836 13240 21864 13280
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 23676 13240 23704 13339
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 24213 13379 24271 13385
rect 24213 13345 24225 13379
rect 24259 13376 24271 13379
rect 24854 13376 24860 13388
rect 24259 13348 24860 13376
rect 24259 13345 24271 13348
rect 24213 13339 24271 13345
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 26970 13336 26976 13388
rect 27028 13376 27034 13388
rect 27065 13379 27123 13385
rect 27065 13376 27077 13379
rect 27028 13348 27077 13376
rect 27028 13336 27034 13348
rect 27065 13345 27077 13348
rect 27111 13345 27123 13379
rect 27065 13339 27123 13345
rect 23753 13311 23811 13317
rect 23753 13277 23765 13311
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 21560 13212 21864 13240
rect 22066 13212 23704 13240
rect 23768 13240 23796 13271
rect 25130 13268 25136 13320
rect 25188 13308 25194 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25188 13280 25237 13308
rect 25188 13268 25194 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 24210 13240 24216 13252
rect 23768 13212 24216 13240
rect 22066 13172 22094 13212
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 18524 13144 22094 13172
rect 23293 13175 23351 13181
rect 23293 13141 23305 13175
rect 23339 13172 23351 13175
rect 23474 13172 23480 13184
rect 23339 13144 23480 13172
rect 23339 13141 23351 13144
rect 23293 13135 23351 13141
rect 23474 13132 23480 13144
rect 23532 13132 23538 13184
rect 1104 13082 28428 13104
rect 1104 13030 5536 13082
rect 5588 13030 5600 13082
rect 5652 13030 5664 13082
rect 5716 13030 5728 13082
rect 5780 13030 14644 13082
rect 14696 13030 14708 13082
rect 14760 13030 14772 13082
rect 14824 13030 14836 13082
rect 14888 13030 23752 13082
rect 23804 13030 23816 13082
rect 23868 13030 23880 13082
rect 23932 13030 23944 13082
rect 23996 13030 28428 13082
rect 1104 13008 28428 13030
rect 4246 12968 4252 12980
rect 4207 12940 4252 12968
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 5644 12940 8217 12968
rect 2774 12792 2780 12844
rect 2832 12832 2838 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2832 12804 2881 12832
rect 2832 12792 2838 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2038 12764 2044 12776
rect 1999 12736 2044 12764
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 3136 12767 3194 12773
rect 3136 12733 3148 12767
rect 3182 12764 3194 12767
rect 4062 12764 4068 12776
rect 3182 12736 4068 12764
rect 3182 12733 3194 12736
rect 3136 12727 3194 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4264 12764 4292 12928
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4264 12736 4721 12764
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 4709 12727 4767 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 5644 12773 5672 12940
rect 8205 12937 8217 12940
rect 8251 12968 8263 12971
rect 8294 12968 8300 12980
rect 8251 12940 8300 12968
rect 8251 12937 8263 12940
rect 8205 12931 8263 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9692 12940 11284 12968
rect 5718 12860 5724 12912
rect 5776 12900 5782 12912
rect 6546 12900 6552 12912
rect 5776 12872 6552 12900
rect 5776 12860 5782 12872
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6696 12804 6837 12832
rect 6696 12792 6702 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 5500 12736 5549 12764
rect 5500 12724 5506 12736
rect 5537 12733 5549 12736
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 5902 12764 5908 12776
rect 5767 12736 5908 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 6656 12764 6684 12792
rect 6420 12736 6684 12764
rect 6420 12724 6426 12736
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8662 12764 8668 12776
rect 8536 12736 8668 12764
rect 8536 12724 8542 12736
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9692 12773 9720 12940
rect 10410 12860 10416 12912
rect 10468 12900 10474 12912
rect 10594 12900 10600 12912
rect 10468 12872 10600 12900
rect 10468 12860 10474 12872
rect 10594 12860 10600 12872
rect 10652 12860 10658 12912
rect 10962 12900 10968 12912
rect 10923 12872 10968 12900
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 11256 12900 11284 12940
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 13906 12968 13912 12980
rect 11388 12940 13912 12968
rect 11388 12928 11394 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 14148 12940 15516 12968
rect 14148 12928 14154 12940
rect 11698 12900 11704 12912
rect 11256 12872 11704 12900
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12250 12900 12256 12912
rect 12124 12872 12256 12900
rect 12124 12860 12130 12872
rect 12250 12860 12256 12872
rect 12308 12900 12314 12912
rect 12308 12872 12434 12900
rect 12308 12860 12314 12872
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 10060 12804 12173 12832
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 7070 12699 7128 12705
rect 7070 12696 7082 12699
rect 5920 12668 7082 12696
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12628 4859 12631
rect 5718 12628 5724 12640
rect 4847 12600 5724 12628
rect 4847 12597 4859 12600
rect 4801 12591 4859 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 5920 12637 5948 12668
rect 7070 12665 7082 12668
rect 7116 12665 7128 12699
rect 7070 12659 7128 12665
rect 7190 12656 7196 12708
rect 7248 12696 7254 12708
rect 7834 12696 7840 12708
rect 7248 12668 7840 12696
rect 7248 12656 7254 12668
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 5905 12631 5963 12637
rect 5905 12597 5917 12631
rect 5951 12597 5963 12631
rect 5905 12591 5963 12597
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6638 12628 6644 12640
rect 6144 12600 6644 12628
rect 6144 12588 6150 12600
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 9508 12628 9536 12727
rect 9784 12696 9812 12727
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10060 12773 10088 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12406 12832 12434 12872
rect 13538 12860 13544 12912
rect 13596 12900 13602 12912
rect 15488 12900 15516 12940
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 15933 12971 15991 12977
rect 15933 12968 15945 12971
rect 15620 12940 15945 12968
rect 15620 12928 15626 12940
rect 15933 12937 15945 12940
rect 15979 12968 15991 12971
rect 18874 12968 18880 12980
rect 15979 12940 18880 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 13596 12872 14596 12900
rect 15488 12872 17540 12900
rect 13596 12860 13602 12872
rect 14568 12832 14596 12872
rect 12406 12804 14412 12832
rect 14568 12804 14688 12832
rect 12161 12795 12219 12801
rect 10045 12767 10103 12773
rect 9916 12736 9961 12764
rect 9916 12724 9922 12736
rect 10045 12733 10057 12767
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 10928 12736 12081 12764
rect 10928 12724 10934 12736
rect 12069 12733 12081 12736
rect 12115 12764 12127 12767
rect 13446 12764 13452 12776
rect 12115 12736 13452 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 14274 12764 14280 12776
rect 13863 12736 14280 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14384 12764 14412 12804
rect 14458 12764 14464 12776
rect 14384 12736 14464 12764
rect 14458 12724 14464 12736
rect 14516 12764 14522 12776
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14516 12736 14565 12764
rect 14516 12724 14522 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 10781 12699 10839 12705
rect 10781 12696 10793 12699
rect 9784 12668 10793 12696
rect 10781 12665 10793 12668
rect 10827 12696 10839 12699
rect 14182 12696 14188 12708
rect 10827 12668 14188 12696
rect 10827 12665 10839 12668
rect 10781 12659 10839 12665
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 6788 12600 9536 12628
rect 6788 12588 6794 12600
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10229 12631 10287 12637
rect 10229 12628 10241 12631
rect 9732 12600 10241 12628
rect 9732 12588 9738 12600
rect 10229 12597 10241 12600
rect 10275 12597 10287 12631
rect 10229 12591 10287 12597
rect 14001 12631 14059 12637
rect 14001 12597 14013 12631
rect 14047 12628 14059 12631
rect 14090 12628 14096 12640
rect 14047 12600 14096 12628
rect 14047 12597 14059 12600
rect 14001 12591 14059 12597
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14660 12628 14688 12804
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 17402 12832 17408 12844
rect 16540 12804 17408 12832
rect 16540 12792 16546 12804
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 17512 12832 17540 12872
rect 17678 12860 17684 12912
rect 17736 12900 17742 12912
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 17736 12872 17785 12900
rect 17736 12860 17742 12872
rect 17773 12869 17785 12872
rect 17819 12900 17831 12903
rect 20254 12900 20260 12912
rect 17819 12872 20260 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 17512 12804 17632 12832
rect 17604 12776 17632 12804
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 21968 12804 23029 12832
rect 21968 12792 21974 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 14820 12767 14878 12773
rect 14820 12733 14832 12767
rect 14866 12764 14878 12767
rect 15286 12764 15292 12776
rect 14866 12736 15292 12764
rect 14866 12733 14878 12736
rect 14820 12727 14878 12733
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 17310 12764 17316 12776
rect 17271 12736 17316 12764
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17497 12767 17555 12773
rect 17497 12733 17509 12767
rect 17543 12733 17555 12767
rect 17497 12727 17555 12733
rect 14918 12656 14924 12708
rect 14976 12696 14982 12708
rect 17512 12696 17540 12727
rect 17586 12724 17592 12776
rect 17644 12764 17650 12776
rect 17865 12767 17923 12773
rect 17644 12736 17737 12764
rect 17644 12724 17650 12736
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18230 12764 18236 12776
rect 17911 12736 18236 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 19610 12764 19616 12776
rect 18380 12736 18425 12764
rect 19571 12736 19616 12764
rect 18380 12724 18386 12736
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19702 12724 19708 12776
rect 19760 12764 19766 12776
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 19760 12736 20269 12764
rect 19760 12724 19766 12736
rect 20257 12733 20269 12736
rect 20303 12733 20315 12767
rect 23032 12764 23060 12795
rect 24946 12764 24952 12776
rect 23032 12736 24952 12764
rect 20257 12727 20315 12733
rect 24946 12724 24952 12736
rect 25004 12764 25010 12776
rect 25130 12764 25136 12776
rect 25004 12736 25136 12764
rect 25004 12724 25010 12736
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 19794 12696 19800 12708
rect 14976 12668 17540 12696
rect 19755 12668 19800 12696
rect 14976 12656 14982 12668
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 20524 12699 20582 12705
rect 20524 12665 20536 12699
rect 20570 12696 20582 12699
rect 20990 12696 20996 12708
rect 20570 12668 20996 12696
rect 20570 12665 20582 12668
rect 20524 12659 20582 12665
rect 20990 12656 20996 12668
rect 21048 12656 21054 12708
rect 23284 12699 23342 12705
rect 23284 12665 23296 12699
rect 23330 12696 23342 12699
rect 23658 12696 23664 12708
rect 23330 12668 23664 12696
rect 23330 12665 23342 12668
rect 23284 12659 23342 12665
rect 23658 12656 23664 12668
rect 23716 12656 23722 12708
rect 25400 12699 25458 12705
rect 25400 12665 25412 12699
rect 25446 12696 25458 12699
rect 25774 12696 25780 12708
rect 25446 12668 25780 12696
rect 25446 12665 25458 12668
rect 25400 12659 25458 12665
rect 25774 12656 25780 12668
rect 25832 12656 25838 12708
rect 16666 12628 16672 12640
rect 14660 12600 16672 12628
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 16816 12600 17325 12628
rect 16816 12588 16822 12600
rect 17313 12597 17325 12600
rect 17359 12597 17371 12631
rect 17313 12591 17371 12597
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 18509 12631 18567 12637
rect 18509 12628 18521 12631
rect 17460 12600 18521 12628
rect 17460 12588 17466 12600
rect 18509 12597 18521 12600
rect 18555 12597 18567 12631
rect 18509 12591 18567 12597
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 20622 12628 20628 12640
rect 20404 12600 20628 12628
rect 20404 12588 20410 12600
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 21634 12628 21640 12640
rect 21595 12600 21640 12628
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 24394 12628 24400 12640
rect 24355 12600 24400 12628
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 25498 12588 25504 12640
rect 25556 12628 25562 12640
rect 26513 12631 26571 12637
rect 26513 12628 26525 12631
rect 25556 12600 26525 12628
rect 25556 12588 25562 12600
rect 26513 12597 26525 12600
rect 26559 12597 26571 12631
rect 26513 12591 26571 12597
rect 1104 12538 28428 12560
rect 1104 12486 10090 12538
rect 10142 12486 10154 12538
rect 10206 12486 10218 12538
rect 10270 12486 10282 12538
rect 10334 12486 19198 12538
rect 19250 12486 19262 12538
rect 19314 12486 19326 12538
rect 19378 12486 19390 12538
rect 19442 12486 28428 12538
rect 1104 12464 28428 12486
rect 8018 12424 8024 12436
rect 6288 12396 8024 12424
rect 2682 12356 2688 12368
rect 1964 12328 2688 12356
rect 1964 12297 1992 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 2216 12291 2274 12297
rect 2216 12257 2228 12291
rect 2262 12288 2274 12291
rect 3694 12288 3700 12300
rect 2262 12260 3700 12288
rect 2262 12257 2274 12260
rect 2216 12251 2274 12257
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4525 12291 4583 12297
rect 4525 12288 4537 12291
rect 4028 12260 4537 12288
rect 4028 12248 4034 12260
rect 4525 12257 4537 12260
rect 4571 12257 4583 12291
rect 4706 12288 4712 12300
rect 4667 12260 4712 12288
rect 4525 12251 4583 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 4890 12288 4896 12300
rect 4851 12260 4896 12288
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6288 12297 6316 12396
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 10686 12424 10692 12436
rect 9784 12396 10692 12424
rect 7193 12359 7251 12365
rect 7193 12325 7205 12359
rect 7239 12356 7251 12359
rect 8570 12356 8576 12368
rect 7239 12328 8576 12356
rect 7239 12325 7251 12328
rect 7193 12319 7251 12325
rect 8570 12316 8576 12328
rect 8628 12316 8634 12368
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6546 12288 6552 12300
rect 6507 12260 6552 12288
rect 6273 12251 6331 12257
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 6104 12220 6132 12251
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 9784 12297 9812 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11698 12424 11704 12436
rect 11659 12396 11704 12424
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 13998 12424 14004 12436
rect 12032 12396 14004 12424
rect 12032 12384 12038 12396
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14918 12424 14924 12436
rect 14879 12396 14924 12424
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 17221 12427 17279 12433
rect 16264 12396 16896 12424
rect 16264 12384 16270 12396
rect 10045 12359 10103 12365
rect 10045 12325 10057 12359
rect 10091 12356 10103 12359
rect 10965 12359 11023 12365
rect 10091 12328 10272 12356
rect 10091 12325 10103 12328
rect 10045 12319 10103 12325
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9950 12288 9956 12300
rect 9863 12260 9956 12288
rect 9769 12251 9827 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10244 12288 10272 12328
rect 10965 12325 10977 12359
rect 11011 12356 11023 12359
rect 11330 12356 11336 12368
rect 11011 12328 11336 12356
rect 11011 12325 11023 12328
rect 10965 12319 11023 12325
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14182 12356 14188 12368
rect 13872 12328 14188 12356
rect 13872 12316 13878 12328
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 15838 12356 15844 12368
rect 15672 12328 15844 12356
rect 10686 12288 10692 12300
rect 10244 12260 10692 12288
rect 10686 12248 10692 12260
rect 10744 12288 10750 12300
rect 11609 12291 11667 12297
rect 11609 12288 11621 12291
rect 10744 12260 11621 12288
rect 10744 12248 10750 12260
rect 11609 12257 11621 12260
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12257 12495 12291
rect 12986 12288 12992 12300
rect 12947 12260 12992 12288
rect 12437 12251 12495 12257
rect 7374 12220 7380 12232
rect 6104 12192 7380 12220
rect 4801 12183 4859 12189
rect 3329 12087 3387 12093
rect 3329 12053 3341 12087
rect 3375 12084 3387 12087
rect 3418 12084 3424 12096
rect 3375 12056 3424 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 4816 12084 4844 12183
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 9968 12220 9996 12248
rect 10778 12220 10784 12232
rect 9968 12192 10784 12220
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 12452 12220 12480 12251
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12288 14887 12291
rect 15010 12288 15016 12300
rect 14875 12260 15016 12288
rect 14875 12257 14887 12260
rect 14829 12251 14887 12257
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 15672 12297 15700 12328
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16022 12288 16028 12300
rect 15804 12260 15849 12288
rect 15983 12260 16028 12288
rect 15804 12248 15810 12260
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16485 12291 16543 12297
rect 16485 12257 16497 12291
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 10928 12192 12480 12220
rect 15473 12223 15531 12229
rect 10928 12180 10934 12192
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 16500 12220 16528 12251
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 16868 12297 16896 12396
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17310 12424 17316 12436
rect 17267 12396 17316 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 18417 12427 18475 12433
rect 18417 12424 18429 12427
rect 18288 12396 18429 12424
rect 18288 12384 18294 12396
rect 18417 12393 18429 12396
rect 18463 12393 18475 12427
rect 18417 12387 18475 12393
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 22005 12427 22063 12433
rect 19852 12396 21956 12424
rect 19852 12384 19858 12396
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 17000 12328 17356 12356
rect 17000 12316 17006 12328
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 16632 12260 16681 12288
rect 16632 12248 16638 12260
rect 16669 12257 16681 12260
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 16853 12291 16911 12297
rect 16853 12257 16865 12291
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 17037 12291 17095 12297
rect 17037 12257 17049 12291
rect 17083 12288 17095 12291
rect 17083 12260 17264 12288
rect 17083 12257 17095 12260
rect 17037 12251 17095 12257
rect 15519 12192 16528 12220
rect 16761 12223 16819 12229
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 16761 12189 16773 12223
rect 16807 12220 16819 12223
rect 16807 12192 16896 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 16868 12164 16896 12192
rect 5261 12155 5319 12161
rect 5261 12121 5273 12155
rect 5307 12152 5319 12155
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5307 12124 5825 12152
rect 5307 12121 5319 12124
rect 5261 12115 5319 12121
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 6365 12155 6423 12161
rect 6365 12152 6377 12155
rect 6328 12124 6377 12152
rect 6328 12112 6334 12124
rect 6365 12121 6377 12124
rect 6411 12121 6423 12155
rect 12066 12152 12072 12164
rect 6365 12115 6423 12121
rect 6472 12124 12072 12152
rect 4982 12084 4988 12096
rect 4816 12056 4988 12084
rect 4982 12044 4988 12056
rect 5040 12084 5046 12096
rect 6472 12084 6500 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 15838 12152 15844 12164
rect 12768 12124 15844 12152
rect 12768 12112 12774 12124
rect 15838 12112 15844 12124
rect 15896 12112 15902 12164
rect 16850 12112 16856 12164
rect 16908 12112 16914 12164
rect 7282 12084 7288 12096
rect 5040 12056 6500 12084
rect 7243 12056 7288 12084
rect 5040 12044 5046 12056
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 10318 12084 10324 12096
rect 10279 12056 10324 12084
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 11054 12084 11060 12096
rect 11015 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 12250 12084 12256 12096
rect 12211 12056 12256 12084
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13354 12084 13360 12096
rect 13127 12056 13360 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 15933 12087 15991 12093
rect 15933 12053 15945 12087
rect 15979 12084 15991 12087
rect 16574 12084 16580 12096
rect 15979 12056 16580 12084
rect 15979 12053 15991 12056
rect 15933 12047 15991 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 17236 12084 17264 12260
rect 17328 12220 17356 12328
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 21266 12356 21272 12368
rect 17644 12328 21272 12356
rect 17644 12316 17650 12328
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 21928 12356 21956 12396
rect 22005 12393 22017 12427
rect 22051 12424 22063 12427
rect 22094 12424 22100 12436
rect 22051 12396 22100 12424
rect 22051 12393 22063 12396
rect 22005 12387 22063 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 22554 12424 22560 12436
rect 22515 12396 22560 12424
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 23474 12424 23480 12436
rect 23308 12396 23480 12424
rect 23308 12365 23336 12396
rect 23474 12384 23480 12396
rect 23532 12384 23538 12436
rect 23658 12424 23664 12436
rect 23619 12396 23664 12424
rect 23658 12384 23664 12396
rect 23716 12384 23722 12436
rect 24210 12424 24216 12436
rect 24171 12396 24216 12424
rect 24210 12384 24216 12396
rect 24268 12384 24274 12436
rect 25774 12424 25780 12436
rect 25735 12396 25780 12424
rect 25774 12384 25780 12396
rect 25832 12384 25838 12436
rect 23293 12359 23351 12365
rect 21928 12328 23152 12356
rect 17678 12288 17684 12300
rect 17639 12260 17684 12288
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 18325 12291 18383 12297
rect 18325 12257 18337 12291
rect 18371 12288 18383 12291
rect 19058 12288 19064 12300
rect 18371 12260 19064 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 19058 12248 19064 12260
rect 19116 12288 19122 12300
rect 20714 12288 20720 12300
rect 19116 12260 20720 12288
rect 19116 12248 19122 12260
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 20892 12291 20950 12297
rect 20892 12257 20904 12291
rect 20938 12288 20950 12291
rect 21174 12288 21180 12300
rect 20938 12260 21180 12288
rect 20938 12257 20950 12260
rect 20892 12251 20950 12257
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 21450 12248 21456 12300
rect 21508 12288 21514 12300
rect 21634 12288 21640 12300
rect 21508 12260 21640 12288
rect 21508 12248 21514 12260
rect 21634 12248 21640 12260
rect 21692 12288 21698 12300
rect 23124 12297 23152 12328
rect 23293 12325 23305 12359
rect 23339 12325 23351 12359
rect 23293 12319 23351 12325
rect 23385 12359 23443 12365
rect 23385 12325 23397 12359
rect 23431 12356 23443 12359
rect 23431 12328 24164 12356
rect 23431 12325 23443 12328
rect 23385 12319 23443 12325
rect 24136 12297 24164 12328
rect 24762 12316 24768 12368
rect 24820 12356 24826 12368
rect 25409 12359 25467 12365
rect 25409 12356 25421 12359
rect 24820 12328 25421 12356
rect 24820 12316 24826 12328
rect 25409 12325 25421 12328
rect 25455 12325 25467 12359
rect 25409 12319 25467 12325
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 26789 12359 26847 12365
rect 26789 12356 26801 12359
rect 26384 12328 26801 12356
rect 26384 12316 26390 12328
rect 26789 12325 26801 12328
rect 26835 12325 26847 12359
rect 26789 12319 26847 12325
rect 26970 12316 26976 12368
rect 27028 12356 27034 12368
rect 27525 12359 27583 12365
rect 27525 12356 27537 12359
rect 27028 12328 27537 12356
rect 27028 12316 27034 12328
rect 27525 12325 27537 12328
rect 27571 12325 27583 12359
rect 27525 12319 27583 12325
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 21692 12260 22477 12288
rect 21692 12248 21698 12260
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22465 12251 22523 12257
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 24121 12291 24179 12297
rect 24121 12257 24133 12291
rect 24167 12288 24179 12291
rect 24394 12288 24400 12300
rect 24167 12260 24400 12288
rect 24167 12257 24179 12260
rect 24121 12251 24179 12257
rect 17586 12220 17592 12232
rect 17328 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 19668 12192 20637 12220
rect 19668 12180 19674 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 23492 12220 23520 12251
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25314 12288 25320 12300
rect 25271 12260 25320 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 25498 12288 25504 12300
rect 25459 12260 25504 12288
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 25593 12291 25651 12297
rect 25593 12257 25605 12291
rect 25639 12257 25651 12291
rect 27706 12288 27712 12300
rect 27667 12260 27712 12288
rect 25593 12251 25651 12257
rect 22704 12192 23520 12220
rect 22704 12180 22710 12192
rect 24210 12180 24216 12232
rect 24268 12220 24274 12232
rect 25608 12220 25636 12251
rect 27706 12248 27712 12260
rect 27764 12248 27770 12300
rect 24268 12192 25636 12220
rect 24268 12180 24274 12192
rect 17773 12155 17831 12161
rect 17773 12121 17785 12155
rect 17819 12152 17831 12155
rect 18690 12152 18696 12164
rect 17819 12124 18696 12152
rect 17819 12121 17831 12124
rect 17773 12115 17831 12121
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 23566 12112 23572 12164
rect 23624 12152 23630 12164
rect 24762 12152 24768 12164
rect 23624 12124 24768 12152
rect 23624 12112 23630 12124
rect 24762 12112 24768 12124
rect 24820 12112 24826 12164
rect 17092 12056 17264 12084
rect 17092 12044 17098 12056
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 25314 12084 25320 12096
rect 18196 12056 25320 12084
rect 18196 12044 18202 12056
rect 25314 12044 25320 12056
rect 25372 12044 25378 12096
rect 26878 12084 26884 12096
rect 26839 12056 26884 12084
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 1104 11994 28428 12016
rect 1104 11942 5536 11994
rect 5588 11942 5600 11994
rect 5652 11942 5664 11994
rect 5716 11942 5728 11994
rect 5780 11942 14644 11994
rect 14696 11942 14708 11994
rect 14760 11942 14772 11994
rect 14824 11942 14836 11994
rect 14888 11942 23752 11994
rect 23804 11942 23816 11994
rect 23868 11942 23880 11994
rect 23932 11942 23944 11994
rect 23996 11942 28428 11994
rect 1104 11920 28428 11942
rect 2746 11852 15792 11880
rect 2222 11772 2228 11824
rect 2280 11812 2286 11824
rect 2746 11812 2774 11852
rect 3694 11812 3700 11824
rect 2280 11784 2774 11812
rect 3655 11784 3700 11812
rect 2280 11772 2286 11784
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 4249 11815 4307 11821
rect 4249 11781 4261 11815
rect 4295 11812 4307 11815
rect 4706 11812 4712 11824
rect 4295 11784 4712 11812
rect 4295 11781 4307 11784
rect 4249 11775 4307 11781
rect 4706 11772 4712 11784
rect 4764 11772 4770 11824
rect 5537 11815 5595 11821
rect 5537 11781 5549 11815
rect 5583 11812 5595 11815
rect 6086 11812 6092 11824
rect 5583 11784 6092 11812
rect 5583 11781 5595 11784
rect 5537 11775 5595 11781
rect 6086 11772 6092 11784
rect 6144 11812 6150 11824
rect 6362 11812 6368 11824
rect 6144 11784 6368 11812
rect 6144 11772 6150 11784
rect 6362 11772 6368 11784
rect 6420 11772 6426 11824
rect 8018 11772 8024 11824
rect 8076 11812 8082 11824
rect 8665 11815 8723 11821
rect 8665 11812 8677 11815
rect 8076 11784 8677 11812
rect 8076 11772 8082 11784
rect 8665 11781 8677 11784
rect 8711 11781 8723 11815
rect 10686 11812 10692 11824
rect 10647 11784 10692 11812
rect 8665 11775 8723 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 12894 11772 12900 11824
rect 12952 11812 12958 11824
rect 13817 11815 13875 11821
rect 12952 11784 13768 11812
rect 12952 11772 12958 11784
rect 9122 11744 9128 11756
rect 1504 11716 9128 11744
rect 1504 11685 1532 11716
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 13354 11744 13360 11756
rect 10428 11716 13032 11744
rect 13315 11716 13360 11744
rect 1489 11679 1547 11685
rect 1489 11645 1501 11679
rect 1535 11645 1547 11679
rect 2130 11676 2136 11688
rect 2091 11648 2136 11676
rect 1489 11639 1547 11645
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 3142 11676 3148 11688
rect 3103 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 3418 11676 3424 11688
rect 3379 11648 3424 11676
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11676 3571 11679
rect 4062 11676 4068 11688
rect 3559 11648 4068 11676
rect 3559 11645 3571 11648
rect 3513 11639 3571 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 5994 11676 6000 11688
rect 5767 11648 6000 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 3329 11611 3387 11617
rect 3329 11608 3341 11611
rect 3292 11580 3341 11608
rect 3292 11568 3298 11580
rect 3329 11577 3341 11580
rect 3375 11577 3387 11611
rect 3436 11608 3464 11636
rect 4172 11608 4200 11639
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11676 6975 11679
rect 8202 11676 8208 11688
rect 6963 11648 8208 11676
rect 6963 11645 6975 11648
rect 6917 11639 6975 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 8812 11648 9321 11676
rect 8812 11636 8818 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9576 11679 9634 11685
rect 9576 11645 9588 11679
rect 9622 11676 9634 11679
rect 10318 11676 10324 11688
rect 9622 11648 10324 11676
rect 9622 11645 9634 11648
rect 9576 11639 9634 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 3436 11580 4200 11608
rect 3329 11571 3387 11577
rect 5350 11568 5356 11620
rect 5408 11608 5414 11620
rect 7282 11608 7288 11620
rect 5408 11580 7288 11608
rect 5408 11568 5414 11580
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 5902 11540 5908 11552
rect 4120 11512 5908 11540
rect 4120 11500 4126 11512
rect 5902 11500 5908 11512
rect 5960 11540 5966 11552
rect 7009 11543 7067 11549
rect 7009 11540 7021 11543
rect 5960 11512 7021 11540
rect 5960 11500 5966 11512
rect 7009 11509 7021 11512
rect 7055 11509 7067 11543
rect 8220 11540 8248 11636
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 10428 11608 10456 11716
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12894 11676 12900 11688
rect 12124 11648 12900 11676
rect 12124 11636 12130 11648
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 8527 11580 10456 11608
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 11974 11608 11980 11620
rect 11388 11580 11980 11608
rect 11388 11568 11394 11580
rect 11974 11568 11980 11580
rect 12032 11568 12038 11620
rect 12161 11611 12219 11617
rect 12161 11577 12173 11611
rect 12207 11577 12219 11611
rect 12161 11571 12219 11577
rect 12345 11611 12403 11617
rect 12345 11577 12357 11611
rect 12391 11608 12403 11611
rect 12618 11608 12624 11620
rect 12391 11580 12624 11608
rect 12391 11577 12403 11580
rect 12345 11571 12403 11577
rect 12176 11540 12204 11571
rect 12618 11568 12624 11580
rect 12676 11568 12682 11620
rect 13004 11608 13032 11716
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13170 11676 13176 11688
rect 13131 11648 13176 11676
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13504 11648 13645 11676
rect 13504 11636 13510 11648
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13740 11676 13768 11784
rect 13817 11781 13829 11815
rect 13863 11812 13875 11815
rect 14734 11812 14740 11824
rect 13863 11784 14740 11812
rect 13863 11781 13875 11784
rect 13817 11775 13875 11781
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 14274 11744 14280 11756
rect 13955 11716 14280 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 15764 11685 15792 11852
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 21174 11880 21180 11892
rect 15896 11852 20668 11880
rect 21135 11852 21180 11880
rect 15896 11840 15902 11852
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 16850 11812 16856 11824
rect 16632 11784 16856 11812
rect 16632 11772 16638 11784
rect 16850 11772 16856 11784
rect 16908 11772 16914 11824
rect 20254 11744 20260 11756
rect 16040 11716 17448 11744
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 13740 11648 14013 11676
rect 13633 11639 13691 11645
rect 14001 11645 14013 11648
rect 14047 11676 14059 11679
rect 15749 11679 15807 11685
rect 14047 11648 15700 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 13814 11608 13820 11620
rect 13004 11580 13820 11608
rect 13814 11568 13820 11580
rect 13872 11608 13878 11620
rect 14090 11608 14096 11620
rect 13872 11580 14096 11608
rect 13872 11568 13878 11580
rect 14090 11568 14096 11580
rect 14148 11568 14154 11620
rect 15672 11608 15700 11648
rect 15749 11645 15761 11679
rect 15795 11645 15807 11679
rect 15930 11676 15936 11688
rect 15891 11648 15936 11676
rect 15749 11639 15807 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16040 11608 16068 11716
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 17126 11676 17132 11688
rect 17000 11648 17132 11676
rect 17000 11636 17006 11648
rect 17126 11636 17132 11648
rect 17184 11676 17190 11688
rect 17313 11679 17371 11685
rect 17313 11676 17325 11679
rect 17184 11648 17325 11676
rect 17184 11636 17190 11648
rect 17313 11645 17325 11648
rect 17359 11645 17371 11679
rect 17420 11676 17448 11716
rect 19444 11716 20260 11744
rect 17954 11676 17960 11688
rect 17420 11648 17960 11676
rect 17313 11639 17371 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 19444 11685 19472 11716
rect 20254 11704 20260 11716
rect 20312 11744 20318 11756
rect 20640 11744 20668 11852
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 24578 11880 24584 11892
rect 21284 11852 24584 11880
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 21284 11812 21312 11852
rect 24578 11840 24584 11852
rect 24636 11840 24642 11892
rect 24854 11880 24860 11892
rect 24815 11852 24860 11880
rect 24854 11840 24860 11852
rect 24912 11840 24918 11892
rect 24946 11840 24952 11892
rect 25004 11880 25010 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 25004 11852 25421 11880
rect 25004 11840 25010 11852
rect 25409 11849 25421 11852
rect 25455 11880 25467 11883
rect 26142 11880 26148 11892
rect 25455 11852 26148 11880
rect 25455 11849 25467 11852
rect 25409 11843 25467 11849
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 20772 11784 21312 11812
rect 21376 11784 26096 11812
rect 20772 11772 20778 11784
rect 21376 11744 21404 11784
rect 20312 11716 20576 11744
rect 20640 11716 21404 11744
rect 20312 11704 20318 11716
rect 19429 11679 19487 11685
rect 19429 11645 19441 11679
rect 19475 11645 19487 11679
rect 20070 11676 20076 11688
rect 20031 11648 20076 11676
rect 19429 11639 19487 11645
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 15672 11580 16068 11608
rect 16117 11611 16175 11617
rect 16117 11577 16129 11611
rect 16163 11608 16175 11611
rect 16574 11608 16580 11620
rect 16163 11580 16580 11608
rect 16163 11577 16175 11580
rect 16117 11571 16175 11577
rect 16574 11568 16580 11580
rect 16632 11568 16638 11620
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 17558 11611 17616 11617
rect 17558 11608 17570 11611
rect 17460 11580 17570 11608
rect 17460 11568 17466 11580
rect 17558 11577 17570 11580
rect 17604 11577 17616 11611
rect 17558 11571 17616 11577
rect 18046 11568 18052 11620
rect 18104 11608 18110 11620
rect 20088 11608 20116 11636
rect 18104 11580 18736 11608
rect 18104 11568 18110 11580
rect 13078 11540 13084 11552
rect 8220 11512 13084 11540
rect 7009 11503 7067 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 18138 11540 18144 11552
rect 13596 11512 18144 11540
rect 13596 11500 13602 11512
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 18708 11549 18736 11580
rect 19260 11580 20116 11608
rect 19260 11549 19288 11580
rect 18693 11543 18751 11549
rect 18693 11509 18705 11543
rect 18739 11509 18751 11543
rect 18693 11503 18751 11509
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11509 19303 11543
rect 19245 11503 19303 11509
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 19668 11512 19901 11540
rect 19668 11500 19674 11512
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 20548 11540 20576 11716
rect 21542 11704 21548 11756
rect 21600 11744 21606 11756
rect 21600 11716 26004 11744
rect 21600 11704 21606 11716
rect 20622 11636 20628 11688
rect 20680 11676 20686 11688
rect 20993 11679 21051 11685
rect 20680 11648 20725 11676
rect 20680 11636 20686 11648
rect 20993 11645 21005 11679
rect 21039 11676 21051 11679
rect 21174 11676 21180 11688
rect 21039 11648 21180 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 23201 11679 23259 11685
rect 23201 11645 23213 11679
rect 23247 11676 23259 11679
rect 23474 11676 23480 11688
rect 23247 11648 23480 11676
rect 23247 11645 23259 11648
rect 23201 11639 23259 11645
rect 23474 11636 23480 11648
rect 23532 11636 23538 11688
rect 24029 11679 24087 11685
rect 24029 11645 24041 11679
rect 24075 11645 24087 11679
rect 24029 11639 24087 11645
rect 24765 11679 24823 11685
rect 24765 11645 24777 11679
rect 24811 11676 24823 11679
rect 25498 11676 25504 11688
rect 24811 11648 25504 11676
rect 24811 11645 24823 11648
rect 24765 11639 24823 11645
rect 20806 11608 20812 11620
rect 20767 11580 20812 11608
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 20901 11611 20959 11617
rect 20901 11577 20913 11611
rect 20947 11608 20959 11611
rect 22094 11608 22100 11620
rect 20947 11580 22100 11608
rect 20947 11577 20959 11580
rect 20901 11571 20959 11577
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 24044 11608 24072 11639
rect 25498 11636 25504 11648
rect 25556 11636 25562 11688
rect 25593 11679 25651 11685
rect 25593 11645 25605 11679
rect 25639 11645 25651 11679
rect 25593 11639 25651 11645
rect 25608 11608 25636 11639
rect 23032 11580 24072 11608
rect 24412 11580 25636 11608
rect 25976 11608 26004 11716
rect 26068 11685 26096 11784
rect 27246 11744 27252 11756
rect 26252 11716 27252 11744
rect 26053 11679 26111 11685
rect 26053 11645 26065 11679
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 26252 11620 26280 11716
rect 27246 11704 27252 11716
rect 27304 11704 27310 11756
rect 26421 11679 26479 11685
rect 26421 11645 26433 11679
rect 26467 11676 26479 11679
rect 26510 11676 26516 11688
rect 26467 11648 26516 11676
rect 26467 11645 26479 11648
rect 26421 11639 26479 11645
rect 26510 11636 26516 11648
rect 26568 11636 26574 11688
rect 26234 11608 26240 11620
rect 25976 11580 26240 11608
rect 23032 11540 23060 11580
rect 24412 11552 24440 11580
rect 26234 11568 26240 11580
rect 26292 11568 26298 11620
rect 26329 11611 26387 11617
rect 26329 11577 26341 11611
rect 26375 11577 26387 11611
rect 26329 11571 26387 11577
rect 23290 11540 23296 11552
rect 20548 11512 23060 11540
rect 23251 11512 23296 11540
rect 19889 11503 19947 11509
rect 23290 11500 23296 11512
rect 23348 11500 23354 11552
rect 23845 11543 23903 11549
rect 23845 11509 23857 11543
rect 23891 11540 23903 11543
rect 24394 11540 24400 11552
rect 23891 11512 24400 11540
rect 23891 11509 23903 11512
rect 23845 11503 23903 11509
rect 24394 11500 24400 11512
rect 24452 11500 24458 11552
rect 25590 11500 25596 11552
rect 25648 11540 25654 11552
rect 26344 11540 26372 11571
rect 26602 11540 26608 11552
rect 25648 11512 26372 11540
rect 26563 11512 26608 11540
rect 25648 11500 25654 11512
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 1104 11450 28428 11472
rect 1104 11398 10090 11450
rect 10142 11398 10154 11450
rect 10206 11398 10218 11450
rect 10270 11398 10282 11450
rect 10334 11398 19198 11450
rect 19250 11398 19262 11450
rect 19314 11398 19326 11450
rect 19378 11398 19390 11450
rect 19442 11398 28428 11450
rect 1104 11376 28428 11398
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 2188 11308 5948 11336
rect 2188 11296 2194 11308
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 5920 11268 5948 11308
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6052 11308 6929 11336
rect 6052 11296 6058 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 13538 11336 13544 11348
rect 8260 11308 13544 11336
rect 8260 11296 8266 11308
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 14274 11336 14280 11348
rect 13771 11308 14280 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15378 11296 15384 11348
rect 15436 11336 15442 11348
rect 15562 11336 15568 11348
rect 15436 11308 15568 11336
rect 15436 11296 15442 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 17402 11336 17408 11348
rect 17359 11308 17408 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17402 11296 17408 11308
rect 17460 11296 17466 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 18012 11308 18245 11336
rect 18012 11296 18018 11308
rect 18233 11305 18245 11308
rect 18279 11336 18291 11339
rect 20622 11336 20628 11348
rect 18279 11308 20628 11336
rect 18279 11305 18291 11308
rect 18233 11299 18291 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 20990 11296 20996 11348
rect 21048 11336 21054 11348
rect 21085 11339 21143 11345
rect 21085 11336 21097 11339
rect 21048 11308 21097 11336
rect 21048 11296 21054 11308
rect 21085 11305 21097 11308
rect 21131 11305 21143 11339
rect 23474 11336 23480 11348
rect 21085 11299 21143 11305
rect 22572 11308 23480 11336
rect 11330 11268 11336 11280
rect 4571 11240 5764 11268
rect 5920 11240 11336 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4430 11200 4436 11212
rect 4391 11172 4436 11200
rect 4249 11163 4307 11169
rect 4264 11132 4292 11163
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5074 11200 5080 11212
rect 4663 11172 5080 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5736 11209 5764 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 11974 11268 11980 11280
rect 11900 11240 11980 11268
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 5902 11200 5908 11212
rect 5767 11172 5908 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8294 11200 8300 11212
rect 8159 11172 8300 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 4338 11132 4344 11144
rect 4264 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 7006 11064 7012 11076
rect 5859 11036 7012 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7116 11064 7144 11163
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 9674 11200 9680 11212
rect 8527 11172 9680 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10312 11203 10370 11209
rect 10312 11169 10324 11203
rect 10358 11200 10370 11203
rect 11146 11200 11152 11212
rect 10358 11172 11152 11200
rect 10358 11169 10370 11172
rect 10312 11163 10370 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11790 11200 11796 11212
rect 11296 11172 11796 11200
rect 11296 11160 11302 11172
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 11900 11209 11928 11240
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 12161 11271 12219 11277
rect 12161 11237 12173 11271
rect 12207 11268 12219 11271
rect 13446 11268 13452 11280
rect 12207 11240 13452 11268
rect 12207 11237 12219 11240
rect 12161 11231 12219 11237
rect 13446 11228 13452 11240
rect 13504 11268 13510 11280
rect 14921 11271 14979 11277
rect 13504 11240 13676 11268
rect 13504 11228 13510 11240
rect 11885 11203 11943 11209
rect 11885 11169 11897 11203
rect 11931 11169 11943 11203
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 11885 11163 11943 11169
rect 11992 11172 12081 11200
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 7432 11104 8401 11132
rect 7432 11092 7438 11104
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 9030 11132 9036 11144
rect 8389 11095 8447 11101
rect 8496 11104 9036 11132
rect 8496 11064 8524 11104
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9950 11132 9956 11144
rect 9180 11104 9956 11132
rect 9180 11092 9186 11104
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 11330 11132 11336 11144
rect 10045 11095 10103 11101
rect 11164 11104 11336 11132
rect 7116 11036 8524 11064
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 10060 11064 10088 11095
rect 11164 11064 11192 11104
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 11992 11132 12020 11172
rect 12069 11169 12081 11172
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 12618 11200 12624 11212
rect 12299 11172 12624 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12894 11200 12900 11212
rect 12855 11172 12900 11200
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 13648 11209 13676 11240
rect 14921 11237 14933 11271
rect 14967 11268 14979 11271
rect 15194 11268 15200 11280
rect 14967 11240 15200 11268
rect 14967 11237 14979 11240
rect 14921 11231 14979 11237
rect 15194 11228 15200 11240
rect 15252 11268 15258 11280
rect 16482 11268 16488 11280
rect 15252 11240 16488 11268
rect 15252 11228 15258 11240
rect 13625 11203 13683 11209
rect 13625 11169 13637 11203
rect 13671 11169 13683 11203
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 13625 11163 13683 11169
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15378 11200 15384 11212
rect 15151 11172 15384 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 14366 11132 14372 11144
rect 11664 11104 12020 11132
rect 12084 11104 14372 11132
rect 11664 11092 11670 11104
rect 8812 11036 10088 11064
rect 8812 11024 8818 11036
rect 4798 10996 4804 11008
rect 4759 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 8205 10999 8263 11005
rect 8205 10965 8217 10999
rect 8251 10996 8263 10999
rect 8478 10996 8484 11008
rect 8251 10968 8484 10996
rect 8251 10965 8263 10968
rect 8205 10959 8263 10965
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 8573 10999 8631 11005
rect 8573 10965 8585 10999
rect 8619 10996 8631 10999
rect 9490 10996 9496 11008
rect 8619 10968 9496 10996
rect 8619 10965 8631 10968
rect 8573 10959 8631 10965
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 10060 10996 10088 11036
rect 10980 11036 11192 11064
rect 10980 10996 11008 11036
rect 11238 11024 11244 11076
rect 11296 11064 11302 11076
rect 11440 11064 11468 11092
rect 12084 11064 12112 11104
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 15028 11132 15056 11163
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15764 11209 15792 11240
rect 16482 11228 16488 11240
rect 16540 11268 16546 11280
rect 16945 11271 17003 11277
rect 16945 11268 16957 11271
rect 16540 11240 16957 11268
rect 16540 11228 16546 11240
rect 16945 11237 16957 11240
rect 16991 11237 17003 11271
rect 16945 11231 17003 11237
rect 17037 11271 17095 11277
rect 17037 11237 17049 11271
rect 17083 11268 17095 11271
rect 19886 11268 19892 11280
rect 17083 11240 19892 11268
rect 17083 11237 17095 11240
rect 17037 11231 17095 11237
rect 19886 11228 19892 11240
rect 19944 11228 19950 11280
rect 20809 11271 20867 11277
rect 20809 11237 20821 11271
rect 20855 11268 20867 11271
rect 21450 11268 21456 11280
rect 20855 11240 21456 11268
rect 20855 11237 20867 11240
rect 20809 11231 20867 11237
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 22186 11228 22192 11280
rect 22244 11268 22250 11280
rect 22572 11277 22600 11308
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 24578 11296 24584 11348
rect 24636 11336 24642 11348
rect 26326 11336 26332 11348
rect 24636 11308 26332 11336
rect 24636 11296 24642 11308
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 26510 11296 26516 11348
rect 26568 11336 26574 11348
rect 27709 11339 27767 11345
rect 27709 11336 27721 11339
rect 26568 11308 27721 11336
rect 26568 11296 26574 11308
rect 27709 11305 27721 11308
rect 27755 11305 27767 11339
rect 27709 11299 27767 11305
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22244 11240 22477 11268
rect 22244 11228 22250 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 22557 11271 22615 11277
rect 22557 11237 22569 11271
rect 22603 11237 22615 11271
rect 22557 11231 22615 11237
rect 23106 11228 23112 11280
rect 23164 11268 23170 11280
rect 23385 11271 23443 11277
rect 23385 11268 23397 11271
rect 23164 11240 23397 11268
rect 23164 11228 23170 11240
rect 23385 11237 23397 11240
rect 23431 11237 23443 11271
rect 25590 11268 25596 11280
rect 25551 11240 25596 11268
rect 23385 11231 23443 11237
rect 25590 11228 25596 11240
rect 25648 11228 25654 11280
rect 26602 11277 26608 11280
rect 26596 11268 26608 11277
rect 26563 11240 26608 11268
rect 26596 11231 26608 11240
rect 26602 11228 26608 11231
rect 26660 11228 26666 11280
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 16758 11200 16764 11212
rect 16719 11172 16764 11200
rect 15749 11163 15807 11169
rect 16758 11160 16764 11172
rect 16816 11160 16822 11212
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 16868 11172 17141 11200
rect 14424 11104 15056 11132
rect 14424 11092 14430 11104
rect 11296 11036 12112 11064
rect 11296 11024 11302 11036
rect 12158 11024 12164 11076
rect 12216 11064 12222 11076
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12216 11036 13093 11064
rect 12216 11024 12222 11036
rect 13081 11033 13093 11036
rect 13127 11033 13139 11067
rect 13081 11027 13139 11033
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13630 11064 13636 11076
rect 13228 11036 13636 11064
rect 13228 11024 13234 11036
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 15102 11064 15108 11076
rect 15015 11036 15108 11064
rect 11422 10996 11428 11008
rect 10060 10968 11008 10996
rect 11383 10968 11428 10996
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12492 10968 12537 10996
rect 12492 10956 12498 10968
rect 12986 10956 12992 11008
rect 13044 10996 13050 11008
rect 15019 10996 15047 11036
rect 15102 11024 15108 11036
rect 15160 11064 15166 11076
rect 15933 11067 15991 11073
rect 15933 11064 15945 11067
rect 15160 11036 15945 11064
rect 15160 11024 15166 11036
rect 15933 11033 15945 11036
rect 15979 11033 15991 11067
rect 15933 11027 15991 11033
rect 15286 10996 15292 11008
rect 13044 10968 15047 10996
rect 15247 10968 15292 10996
rect 13044 10956 13050 10968
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 15948 10996 15976 11027
rect 16022 11024 16028 11076
rect 16080 11064 16086 11076
rect 16666 11064 16672 11076
rect 16080 11036 16672 11064
rect 16080 11024 16086 11036
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 16758 11024 16764 11076
rect 16816 11064 16822 11076
rect 16868 11064 16896 11172
rect 17129 11169 17141 11172
rect 17175 11200 17187 11203
rect 17954 11200 17960 11212
rect 17175 11172 17960 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18414 11200 18420 11212
rect 18095 11172 18420 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 20438 11200 20444 11212
rect 18923 11172 20444 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 20533 11203 20591 11209
rect 20533 11169 20545 11203
rect 20579 11169 20591 11203
rect 20714 11200 20720 11212
rect 20675 11172 20720 11200
rect 20533 11163 20591 11169
rect 16816 11036 16896 11064
rect 16960 11104 19748 11132
rect 16816 11024 16822 11036
rect 16960 10996 16988 11104
rect 17126 11024 17132 11076
rect 17184 11064 17190 11076
rect 19610 11064 19616 11076
rect 17184 11036 19616 11064
rect 17184 11024 17190 11036
rect 19610 11024 19616 11036
rect 19668 11024 19674 11076
rect 19720 11064 19748 11104
rect 19794 11092 19800 11144
rect 19852 11132 19858 11144
rect 20548 11132 20576 11163
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 22281 11203 22339 11209
rect 22281 11200 22293 11203
rect 22066 11172 22293 11200
rect 22066 11132 22094 11172
rect 22281 11169 22293 11172
rect 22327 11169 22339 11203
rect 22646 11200 22652 11212
rect 22281 11163 22339 11169
rect 22388 11172 22652 11200
rect 19852 11104 22094 11132
rect 19852 11092 19858 11104
rect 21542 11064 21548 11076
rect 19720 11036 21548 11064
rect 21542 11024 21548 11036
rect 21600 11024 21606 11076
rect 15948 10968 16988 10996
rect 17402 10956 17408 11008
rect 17460 10996 17466 11008
rect 17586 10996 17592 11008
rect 17460 10968 17592 10996
rect 17460 10956 17466 10968
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 18414 10956 18420 11008
rect 18472 10996 18478 11008
rect 18969 10999 19027 11005
rect 18969 10996 18981 10999
rect 18472 10968 18981 10996
rect 18472 10956 18478 10968
rect 18969 10965 18981 10968
rect 19015 10965 19027 10999
rect 18969 10959 19027 10965
rect 20898 10956 20904 11008
rect 20956 10996 20962 11008
rect 21910 10996 21916 11008
rect 20956 10968 21916 10996
rect 20956 10956 20962 10968
rect 21910 10956 21916 10968
rect 21968 10996 21974 11008
rect 22388 10996 22416 11172
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11169 23351 11203
rect 23750 11200 23756 11212
rect 23711 11172 23756 11200
rect 23293 11163 23351 11169
rect 22738 11024 22744 11076
rect 22796 11064 22802 11076
rect 23014 11064 23020 11076
rect 22796 11036 23020 11064
rect 22796 11024 22802 11036
rect 23014 11024 23020 11036
rect 23072 11024 23078 11076
rect 23308 11064 23336 11163
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 24118 11200 24124 11212
rect 24079 11172 24124 11200
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 24305 11203 24363 11209
rect 24305 11169 24317 11203
rect 24351 11200 24363 11203
rect 24946 11200 24952 11212
rect 24351 11172 24952 11200
rect 24351 11169 24363 11172
rect 24305 11163 24363 11169
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 25314 11200 25320 11212
rect 25275 11172 25320 11200
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 25501 11203 25559 11209
rect 25501 11169 25513 11203
rect 25547 11169 25559 11203
rect 25682 11200 25688 11212
rect 25643 11172 25688 11200
rect 25501 11163 25559 11169
rect 23845 11135 23903 11141
rect 23845 11101 23857 11135
rect 23891 11132 23903 11135
rect 24210 11132 24216 11144
rect 23891 11104 24216 11132
rect 23891 11101 23903 11104
rect 23845 11095 23903 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 25516 11132 25544 11163
rect 25682 11160 25688 11172
rect 25740 11160 25746 11212
rect 26142 11160 26148 11212
rect 26200 11200 26206 11212
rect 26329 11203 26387 11209
rect 26329 11200 26341 11203
rect 26200 11172 26341 11200
rect 26200 11160 26206 11172
rect 26329 11169 26341 11172
rect 26375 11169 26387 11203
rect 26329 11163 26387 11169
rect 26234 11132 26240 11144
rect 25516 11104 26240 11132
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 24302 11064 24308 11076
rect 23308 11036 24308 11064
rect 24302 11024 24308 11036
rect 24360 11024 24366 11076
rect 22830 10996 22836 11008
rect 21968 10968 22416 10996
rect 22791 10968 22836 10996
rect 21968 10956 21974 10968
rect 22830 10956 22836 10968
rect 22888 10956 22894 11008
rect 25774 10956 25780 11008
rect 25832 10996 25838 11008
rect 25869 10999 25927 11005
rect 25869 10996 25881 10999
rect 25832 10968 25881 10996
rect 25832 10956 25838 10968
rect 25869 10965 25881 10968
rect 25915 10965 25927 10999
rect 25869 10959 25927 10965
rect 1104 10906 28428 10928
rect 1104 10854 5536 10906
rect 5588 10854 5600 10906
rect 5652 10854 5664 10906
rect 5716 10854 5728 10906
rect 5780 10854 14644 10906
rect 14696 10854 14708 10906
rect 14760 10854 14772 10906
rect 14824 10854 14836 10906
rect 14888 10854 23752 10906
rect 23804 10854 23816 10906
rect 23868 10854 23880 10906
rect 23932 10854 23944 10906
rect 23996 10854 28428 10906
rect 1104 10832 28428 10854
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10008 10764 10149 10792
rect 10008 10752 10014 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 11146 10792 11152 10804
rect 11107 10764 11152 10792
rect 10137 10755 10195 10761
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 12342 10792 12348 10804
rect 12084 10764 12348 10792
rect 4890 10684 4896 10736
rect 4948 10724 4954 10736
rect 4948 10696 5120 10724
rect 4948 10684 4954 10696
rect 1670 10616 1676 10668
rect 1728 10656 1734 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 1728 10628 2697 10656
rect 1728 10616 1734 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 4982 10656 4988 10668
rect 4943 10628 4988 10656
rect 2685 10619 2743 10625
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2130 10588 2136 10600
rect 1903 10560 2136 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 2700 10588 2728 10619
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5092 10665 5120 10696
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 8297 10727 8355 10733
rect 8297 10724 8309 10727
rect 8260 10696 8309 10724
rect 8260 10684 8266 10696
rect 8297 10693 8309 10696
rect 8343 10693 8355 10727
rect 8297 10687 8355 10693
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 12084 10724 12112 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13446 10792 13452 10804
rect 13407 10764 13452 10792
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 16114 10792 16120 10804
rect 13964 10764 16120 10792
rect 13964 10752 13970 10764
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 24946 10792 24952 10804
rect 24907 10764 24952 10792
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 11388 10696 12112 10724
rect 11388 10684 11394 10696
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 7006 10656 7012 10668
rect 6967 10628 7012 10656
rect 5077 10619 5135 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 8018 10656 8024 10668
rect 7300 10628 8024 10656
rect 3510 10588 3516 10600
rect 2700 10560 3516 10588
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 4706 10588 4712 10600
rect 4667 10560 4712 10588
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4890 10588 4896 10600
rect 4851 10560 4896 10588
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5258 10588 5264 10600
rect 5219 10560 5264 10588
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 7300 10597 7328 10628
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8754 10656 8760 10668
rect 8715 10628 8760 10656
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 11054 10656 11060 10668
rect 10612 10628 11060 10656
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 10612 10597 10640 10628
rect 11054 10616 11060 10628
rect 11112 10656 11118 10668
rect 11974 10656 11980 10668
rect 11112 10628 11980 10656
rect 11112 10616 11118 10628
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12084 10665 12112 10696
rect 16206 10684 16212 10736
rect 16264 10724 16270 10736
rect 16942 10724 16948 10736
rect 16264 10696 16948 10724
rect 16264 10684 16270 10696
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 17586 10684 17592 10736
rect 17644 10724 17650 10736
rect 17862 10724 17868 10736
rect 17644 10696 17868 10724
rect 17644 10684 17650 10696
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14516 10628 14657 10656
rect 14516 10616 14522 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 17368 10628 18153 10656
rect 17368 10616 17374 10628
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 18141 10619 18199 10625
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18506 10656 18512 10668
rect 18279 10628 18512 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 19610 10656 19616 10668
rect 19571 10628 19616 10656
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7432 10560 7573 10588
rect 7432 10548 7438 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 10778 10588 10784 10600
rect 10739 10560 10784 10588
rect 10597 10551 10655 10557
rect 2952 10523 3010 10529
rect 2952 10489 2964 10523
rect 2998 10520 3010 10523
rect 4522 10520 4528 10532
rect 2998 10492 4528 10520
rect 2998 10489 3010 10492
rect 2952 10483 3010 10489
rect 4522 10480 4528 10492
rect 4580 10480 4586 10532
rect 5445 10523 5503 10529
rect 5445 10489 5457 10523
rect 5491 10520 5503 10523
rect 7944 10520 7972 10551
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 14912 10591 14970 10597
rect 11011 10560 11744 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 5491 10492 7972 10520
rect 9024 10523 9082 10529
rect 5491 10489 5503 10492
rect 5445 10483 5503 10489
rect 9024 10489 9036 10523
rect 9070 10520 9082 10523
rect 9950 10520 9956 10532
rect 9070 10492 9956 10520
rect 9070 10489 9082 10492
rect 9024 10483 9082 10489
rect 9950 10480 9956 10492
rect 10008 10480 10014 10532
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10520 10931 10523
rect 11422 10520 11428 10532
rect 10919 10492 11428 10520
rect 10919 10489 10931 10492
rect 10873 10483 10931 10489
rect 11422 10480 11428 10492
rect 11480 10480 11486 10532
rect 1946 10452 1952 10464
rect 1907 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4246 10452 4252 10464
rect 4111 10424 4252 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 11716 10452 11744 10560
rect 14912 10557 14924 10591
rect 14958 10588 14970 10591
rect 15286 10588 15292 10600
rect 14958 10560 15292 10588
rect 14958 10557 14970 10560
rect 14912 10551 14970 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 17862 10588 17868 10600
rect 17823 10560 17868 10588
rect 17862 10548 17868 10560
rect 17920 10548 17926 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18049 10551 18107 10557
rect 12336 10523 12394 10529
rect 12336 10489 12348 10523
rect 12382 10520 12394 10523
rect 12434 10520 12440 10532
rect 12382 10492 12440 10520
rect 12382 10489 12394 10492
rect 12336 10483 12394 10489
rect 12434 10480 12440 10492
rect 12492 10480 12498 10532
rect 14001 10523 14059 10529
rect 14001 10489 14013 10523
rect 14047 10520 14059 10523
rect 15194 10520 15200 10532
rect 14047 10492 15200 10520
rect 14047 10489 14059 10492
rect 14001 10483 14059 10489
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 18064 10520 18092 10551
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 22741 10591 22799 10597
rect 22741 10557 22753 10591
rect 22787 10588 22799 10591
rect 24857 10591 24915 10597
rect 22787 10560 22968 10588
rect 22787 10557 22799 10560
rect 22741 10551 22799 10557
rect 18708 10520 18736 10548
rect 18064 10492 18736 10520
rect 19880 10523 19938 10529
rect 19880 10489 19892 10523
rect 19926 10520 19938 10523
rect 20714 10520 20720 10532
rect 19926 10492 20720 10520
rect 19926 10489 19938 10492
rect 19880 10483 19938 10489
rect 20714 10480 20720 10492
rect 20772 10480 20778 10532
rect 22940 10464 22968 10560
rect 24857 10557 24869 10591
rect 24903 10557 24915 10591
rect 25498 10588 25504 10600
rect 25459 10560 25504 10588
rect 24857 10551 24915 10557
rect 23008 10523 23066 10529
rect 23008 10489 23020 10523
rect 23054 10520 23066 10523
rect 23198 10520 23204 10532
rect 23054 10492 23204 10520
rect 23054 10489 23066 10492
rect 23008 10483 23066 10489
rect 23198 10480 23204 10492
rect 23256 10480 23262 10532
rect 24872 10520 24900 10551
rect 25498 10548 25504 10560
rect 25556 10548 25562 10600
rect 25774 10597 25780 10600
rect 25768 10588 25780 10597
rect 25735 10560 25780 10588
rect 25768 10551 25780 10560
rect 25774 10548 25780 10551
rect 25832 10548 25838 10600
rect 26142 10520 26148 10532
rect 24872 10492 26148 10520
rect 26142 10480 26148 10492
rect 26200 10480 26206 10532
rect 12618 10452 12624 10464
rect 11716 10424 12624 10452
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 13596 10424 14105 10452
rect 13596 10412 13602 10424
rect 14093 10421 14105 10424
rect 14139 10421 14151 10455
rect 14093 10415 14151 10421
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 16025 10455 16083 10461
rect 16025 10452 16037 10455
rect 15436 10424 16037 10452
rect 15436 10412 15442 10424
rect 16025 10421 16037 10424
rect 16071 10452 16083 10455
rect 16114 10452 16120 10464
rect 16071 10424 16120 10452
rect 16071 10421 16083 10424
rect 16025 10415 16083 10421
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 18601 10455 18659 10461
rect 18601 10421 18613 10455
rect 18647 10452 18659 10455
rect 18690 10452 18696 10464
rect 18647 10424 18696 10452
rect 18647 10421 18659 10424
rect 18601 10415 18659 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 20990 10452 20996 10464
rect 20951 10424 20996 10452
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 24118 10452 24124 10464
rect 24079 10424 24124 10452
rect 24118 10412 24124 10424
rect 24176 10412 24182 10464
rect 25682 10412 25688 10464
rect 25740 10452 25746 10464
rect 26881 10455 26939 10461
rect 26881 10452 26893 10455
rect 25740 10424 26893 10452
rect 25740 10412 25746 10424
rect 26881 10421 26893 10424
rect 26927 10421 26939 10455
rect 26881 10415 26939 10421
rect 1104 10362 28428 10384
rect 1104 10310 10090 10362
rect 10142 10310 10154 10362
rect 10206 10310 10218 10362
rect 10270 10310 10282 10362
rect 10334 10310 19198 10362
rect 19250 10310 19262 10362
rect 19314 10310 19326 10362
rect 19378 10310 19390 10362
rect 19442 10310 28428 10362
rect 1104 10288 28428 10310
rect 2866 10248 2872 10260
rect 2827 10220 2872 10248
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5902 10248 5908 10260
rect 5675 10220 5908 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 10008 10220 10057 10248
rect 10008 10208 10014 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10045 10211 10103 10217
rect 17589 10251 17647 10257
rect 17589 10217 17601 10251
rect 17635 10248 17647 10251
rect 17678 10248 17684 10260
rect 17635 10220 17684 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 17920 10220 18153 10248
rect 17920 10208 17926 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 20438 10208 20444 10260
rect 20496 10248 20502 10260
rect 21361 10251 21419 10257
rect 21361 10248 21373 10251
rect 20496 10220 21373 10248
rect 20496 10208 20502 10220
rect 21361 10217 21373 10220
rect 21407 10217 21419 10251
rect 21361 10211 21419 10217
rect 23474 10208 23480 10260
rect 23532 10248 23538 10260
rect 23661 10251 23719 10257
rect 23661 10248 23673 10251
rect 23532 10220 23673 10248
rect 23532 10208 23538 10220
rect 23661 10217 23673 10220
rect 23707 10217 23719 10251
rect 24210 10248 24216 10260
rect 24171 10220 24216 10248
rect 23661 10211 23719 10217
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 26142 10208 26148 10260
rect 26200 10248 26206 10260
rect 26697 10251 26755 10257
rect 26697 10248 26709 10251
rect 26200 10220 26709 10248
rect 26200 10208 26206 10220
rect 26697 10217 26709 10220
rect 26743 10217 26755 10251
rect 26697 10211 26755 10217
rect 4516 10183 4574 10189
rect 4516 10149 4528 10183
rect 4562 10180 4574 10183
rect 4798 10180 4804 10192
rect 4562 10152 4804 10180
rect 4562 10149 4574 10152
rect 4516 10143 4574 10149
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 10597 10183 10655 10189
rect 10597 10180 10609 10183
rect 8352 10152 10609 10180
rect 8352 10140 8358 10152
rect 10597 10149 10609 10152
rect 10643 10149 10655 10183
rect 10597 10143 10655 10149
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12069 10183 12127 10189
rect 12069 10180 12081 10183
rect 12032 10152 12081 10180
rect 12032 10140 12038 10152
rect 12069 10149 12081 10152
rect 12115 10180 12127 10183
rect 12526 10180 12532 10192
rect 12115 10152 12532 10180
rect 12115 10149 12127 10152
rect 12069 10143 12127 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 17126 10180 17132 10192
rect 16224 10152 17132 10180
rect 1756 10115 1814 10121
rect 1756 10081 1768 10115
rect 1802 10112 1814 10115
rect 2682 10112 2688 10124
rect 1802 10084 2688 10112
rect 1802 10081 1814 10084
rect 1756 10075 1814 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3568 10084 4261 10112
rect 3568 10072 3574 10084
rect 4249 10081 4261 10084
rect 4295 10112 4307 10115
rect 4982 10112 4988 10124
rect 4295 10084 4988 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6345 10115 6403 10121
rect 6345 10112 6357 10115
rect 5960 10084 6357 10112
rect 5960 10072 5966 10084
rect 6345 10081 6357 10084
rect 6391 10081 6403 10115
rect 9490 10112 9496 10124
rect 9451 10084 9496 10112
rect 6345 10075 6403 10081
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 9907 10115 9965 10121
rect 9824 10084 9869 10112
rect 9824 10072 9830 10084
rect 9907 10081 9919 10115
rect 9953 10081 9965 10115
rect 9907 10075 9965 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 11422 10112 11428 10124
rect 10551 10084 11428 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10013 1547 10047
rect 6086 10044 6092 10056
rect 6047 10016 6092 10044
rect 1489 10007 1547 10013
rect 1504 9908 1532 10007
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 7926 10044 7932 10056
rect 7616 10016 7932 10044
rect 7616 10004 7622 10016
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9922 10044 9950 10075
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11848 10084 11897 10112
rect 11848 10072 11854 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 12158 10112 12164 10124
rect 12119 10084 12164 10112
rect 11885 10075 11943 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 16224 10121 16252 10152
rect 17126 10140 17132 10152
rect 17184 10140 17190 10192
rect 22548 10183 22606 10189
rect 19996 10152 22094 10180
rect 16209 10115 16267 10121
rect 12308 10084 12353 10112
rect 12308 10072 12314 10084
rect 16209 10081 16221 10115
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 16476 10115 16534 10121
rect 16476 10081 16488 10115
rect 16522 10112 16534 10115
rect 17310 10112 17316 10124
rect 16522 10084 17316 10112
rect 16522 10081 16534 10084
rect 16476 10075 16534 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10081 18383 10115
rect 18325 10075 18383 10081
rect 11238 10044 11244 10056
rect 9922 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 18340 10044 18368 10075
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18693 10115 18751 10121
rect 18472 10084 18517 10112
rect 18472 10072 18478 10084
rect 18693 10081 18705 10115
rect 18739 10112 18751 10115
rect 18874 10112 18880 10124
rect 18739 10084 18880 10112
rect 18739 10081 18751 10084
rect 18693 10075 18751 10081
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19996 10121 20024 10152
rect 19981 10115 20039 10121
rect 19981 10081 19993 10115
rect 20027 10081 20039 10115
rect 19981 10075 20039 10081
rect 20248 10115 20306 10121
rect 20248 10081 20260 10115
rect 20294 10112 20306 10115
rect 20530 10112 20536 10124
rect 20294 10084 20536 10112
rect 20294 10081 20306 10084
rect 20248 10075 20306 10081
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 22066 10112 22094 10152
rect 22548 10149 22560 10183
rect 22594 10180 22606 10183
rect 22830 10180 22836 10192
rect 22594 10152 22836 10180
rect 22594 10149 22606 10152
rect 22548 10143 22606 10149
rect 22830 10140 22836 10152
rect 22888 10140 22894 10192
rect 22922 10140 22928 10192
rect 22980 10180 22986 10192
rect 25498 10180 25504 10192
rect 22980 10152 25504 10180
rect 22980 10140 22986 10152
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 27522 10180 27528 10192
rect 27483 10152 27528 10180
rect 27522 10140 27528 10152
rect 27580 10140 27586 10192
rect 27709 10183 27767 10189
rect 27709 10149 27721 10183
rect 27755 10180 27767 10183
rect 27798 10180 27804 10192
rect 27755 10152 27804 10180
rect 27755 10149 27767 10152
rect 27709 10143 27767 10149
rect 27798 10140 27804 10152
rect 27856 10140 27862 10192
rect 22281 10115 22339 10121
rect 22281 10112 22293 10115
rect 22066 10084 22293 10112
rect 22281 10081 22293 10084
rect 22327 10112 22339 10115
rect 22940 10112 22968 10140
rect 22327 10084 22968 10112
rect 22327 10081 22339 10084
rect 22281 10075 22339 10081
rect 23566 10072 23572 10124
rect 23624 10112 23630 10124
rect 24118 10112 24124 10124
rect 23624 10084 24124 10112
rect 23624 10072 23630 10084
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 25317 10115 25375 10121
rect 25317 10081 25329 10115
rect 25363 10112 25375 10115
rect 25516 10112 25544 10140
rect 25590 10121 25596 10124
rect 25363 10084 25544 10112
rect 25363 10081 25375 10084
rect 25317 10075 25375 10081
rect 25584 10075 25596 10121
rect 25648 10112 25654 10124
rect 25648 10084 25684 10112
rect 25590 10072 25596 10075
rect 25648 10072 25654 10084
rect 19886 10044 19892 10056
rect 18340 10016 19892 10044
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 10318 9936 10324 9988
rect 10376 9976 10382 9988
rect 11606 9976 11612 9988
rect 10376 9948 11612 9976
rect 10376 9936 10382 9948
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12250 9976 12256 9988
rect 11756 9948 12256 9976
rect 11756 9936 11762 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 1670 9908 1676 9920
rect 1504 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 7558 9908 7564 9920
rect 7515 9880 7564 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12526 9908 12532 9920
rect 12483 9880 12532 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 18601 9911 18659 9917
rect 18601 9908 18613 9911
rect 17644 9880 18613 9908
rect 17644 9868 17650 9880
rect 18601 9877 18613 9880
rect 18647 9877 18659 9911
rect 18601 9871 18659 9877
rect 1104 9818 28428 9840
rect 1104 9766 5536 9818
rect 5588 9766 5600 9818
rect 5652 9766 5664 9818
rect 5716 9766 5728 9818
rect 5780 9766 14644 9818
rect 14696 9766 14708 9818
rect 14760 9766 14772 9818
rect 14824 9766 14836 9818
rect 14888 9766 23752 9818
rect 23804 9766 23816 9818
rect 23868 9766 23880 9818
rect 23932 9766 23944 9818
rect 23996 9766 28428 9818
rect 1104 9744 28428 9766
rect 5902 9704 5908 9716
rect 5863 9676 5908 9704
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 20622 9664 20628 9716
rect 20680 9704 20686 9716
rect 20680 9676 20852 9704
rect 20680 9664 20686 9676
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 3200 9608 4476 9636
rect 3200 9596 3206 9608
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 2041 9571 2099 9577
rect 2041 9568 2053 9571
rect 1728 9540 2053 9568
rect 1728 9528 1734 9540
rect 2041 9537 2053 9540
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 3988 9509 4016 9608
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4448 9568 4476 9608
rect 4982 9596 4988 9648
rect 5040 9636 5046 9648
rect 5040 9608 5948 9636
rect 5040 9596 5046 9608
rect 5920 9568 5948 9608
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 10045 9639 10103 9645
rect 10045 9636 10057 9639
rect 10008 9608 10057 9636
rect 10008 9596 10014 9608
rect 10045 9605 10057 9608
rect 10091 9636 10103 9639
rect 10870 9636 10876 9648
rect 10091 9608 10876 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 13817 9639 13875 9645
rect 13817 9605 13829 9639
rect 13863 9636 13875 9639
rect 13906 9636 13912 9648
rect 13863 9608 13912 9636
rect 13863 9605 13875 9608
rect 13817 9599 13875 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 17310 9636 17316 9648
rect 17271 9608 17316 9636
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 19245 9639 19303 9645
rect 17420 9608 19196 9636
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 4120 9540 4384 9568
rect 4448 9540 5396 9568
rect 4120 9528 4126 9540
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 4246 9500 4252 9512
rect 4207 9472 4252 9500
rect 3973 9463 4031 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4356 9509 4384 9540
rect 5368 9512 5396 9540
rect 5644 9540 5856 9568
rect 5920 9540 6837 9568
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 5350 9500 5356 9512
rect 4387 9472 5212 9500
rect 5311 9472 5356 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 2308 9435 2366 9441
rect 2308 9401 2320 9435
rect 2354 9432 2366 9435
rect 2866 9432 2872 9444
rect 2354 9404 2872 9432
rect 2354 9401 2366 9404
rect 2308 9395 2366 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 4157 9435 4215 9441
rect 4157 9432 4169 9435
rect 3344 9404 4169 9432
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2498 9364 2504 9376
rect 1627 9336 2504 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2498 9324 2504 9336
rect 2556 9364 2562 9376
rect 3344 9364 3372 9404
rect 4157 9401 4169 9404
rect 4203 9432 4215 9435
rect 4430 9432 4436 9444
rect 4203 9404 4436 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 2556 9336 3372 9364
rect 3421 9367 3479 9373
rect 2556 9324 2562 9336
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 3602 9364 3608 9376
rect 3467 9336 3608 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 4522 9364 4528 9376
rect 4483 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 5184 9364 5212 9472
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5644 9509 5672 9540
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9469 5779 9503
rect 5828 9500 5856 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 8128 9540 12296 9568
rect 7558 9500 7564 9512
rect 5828 9472 7564 9500
rect 5721 9463 5779 9469
rect 5534 9432 5540 9444
rect 5495 9404 5540 9432
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 5736 9432 5764 9463
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 6730 9432 6736 9444
rect 5736 9404 6736 9432
rect 5736 9364 5764 9404
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6972 9404 7082 9432
rect 6972 9392 6978 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 7070 9395 7128 9401
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 8128 9432 8156 9540
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 7524 9404 8156 9432
rect 8220 9472 8677 9500
rect 7524 9392 7530 9404
rect 5184 9336 5764 9364
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 8220 9373 8248 9472
rect 8665 9469 8677 9472
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 9398 9500 9404 9512
rect 9355 9472 9404 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 10686 9500 10692 9512
rect 10275 9472 10692 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 12158 9500 12164 9512
rect 11011 9472 12164 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 6696 9336 8217 9364
rect 6696 9324 6702 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8754 9364 8760 9376
rect 8715 9336 8760 9364
rect 8205 9327 8263 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 11054 9364 11060 9376
rect 11015 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 12268 9364 12296 9540
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12492 9540 12537 9568
rect 12492 9528 12498 9540
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 17420 9568 17448 9608
rect 13504 9540 17448 9568
rect 13504 9528 13510 9540
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17828 9540 17877 9568
rect 17828 9528 17834 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 12693 9503 12751 9509
rect 12693 9500 12705 9503
rect 12584 9472 12705 9500
rect 12584 9460 12590 9472
rect 12693 9469 12705 9472
rect 12739 9469 12751 9503
rect 12693 9463 12751 9469
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14424 9472 14473 9500
rect 14424 9460 14430 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17310 9500 17316 9512
rect 17000 9472 17316 9500
rect 17000 9460 17006 9472
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 17678 9460 17684 9512
rect 17736 9500 17742 9512
rect 18690 9500 18696 9512
rect 17736 9472 17816 9500
rect 18651 9472 18696 9500
rect 17736 9460 17742 9472
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 14645 9435 14703 9441
rect 14645 9432 14657 9435
rect 13688 9404 14657 9432
rect 13688 9392 13694 9404
rect 14645 9401 14657 9404
rect 14691 9432 14703 9435
rect 15010 9432 15016 9444
rect 14691 9404 15016 9432
rect 14691 9401 14703 9404
rect 14645 9395 14703 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 17788 9441 17816 9472
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 18966 9500 18972 9512
rect 18927 9472 18972 9500
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19168 9509 19196 9608
rect 19245 9605 19257 9639
rect 19291 9636 19303 9639
rect 19518 9636 19524 9648
rect 19291 9608 19524 9636
rect 19291 9605 19303 9608
rect 19245 9599 19303 9605
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 19702 9636 19708 9648
rect 19628 9608 19708 9636
rect 19153 9503 19211 9509
rect 19153 9469 19165 9503
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9500 19579 9503
rect 19628 9500 19656 9608
rect 19702 9596 19708 9608
rect 19760 9636 19766 9648
rect 20254 9636 20260 9648
rect 19760 9608 20260 9636
rect 19760 9596 19766 9608
rect 20254 9596 20260 9608
rect 20312 9596 20318 9648
rect 20714 9636 20720 9648
rect 20675 9608 20720 9636
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 20824 9636 20852 9676
rect 20824 9608 23796 9636
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 21269 9571 21327 9577
rect 21269 9568 21281 9571
rect 19944 9540 21281 9568
rect 19944 9528 19950 9540
rect 21269 9537 21281 9540
rect 21315 9537 21327 9571
rect 23014 9568 23020 9580
rect 22975 9540 23020 9568
rect 21269 9531 21327 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 23290 9568 23296 9580
rect 23251 9540 23296 9568
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 19567 9472 19656 9500
rect 19705 9503 19763 9509
rect 19567 9469 19579 9472
rect 19521 9463 19579 9469
rect 19705 9469 19717 9503
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 20165 9503 20223 9509
rect 20165 9469 20177 9503
rect 20211 9500 20223 9503
rect 20254 9500 20260 9512
rect 20211 9472 20260 9500
rect 20211 9469 20223 9472
rect 20165 9463 20223 9469
rect 17773 9435 17831 9441
rect 17773 9401 17785 9435
rect 17819 9401 17831 9435
rect 17773 9395 17831 9401
rect 13722 9364 13728 9376
rect 12268 9336 13728 9364
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 17678 9364 17684 9376
rect 17639 9336 17684 9364
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 19720 9364 19748 9463
rect 20254 9460 20260 9472
rect 20312 9460 20318 9512
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9500 20591 9503
rect 20898 9500 20904 9512
rect 20579 9472 20904 9500
rect 20579 9469 20591 9472
rect 20533 9463 20591 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 20990 9460 20996 9512
rect 21048 9500 21054 9512
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 21048 9472 21189 9500
rect 21048 9460 21054 9472
rect 21177 9469 21189 9472
rect 21223 9469 21235 9503
rect 22922 9500 22928 9512
rect 22883 9472 22928 9500
rect 21177 9463 21235 9469
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23106 9460 23112 9512
rect 23164 9500 23170 9512
rect 23768 9509 23796 9608
rect 23385 9503 23443 9509
rect 23385 9500 23397 9503
rect 23164 9472 23397 9500
rect 23164 9460 23170 9472
rect 23385 9469 23397 9472
rect 23431 9469 23443 9503
rect 23385 9463 23443 9469
rect 23753 9503 23811 9509
rect 23753 9469 23765 9503
rect 23799 9469 23811 9503
rect 23753 9463 23811 9469
rect 23937 9503 23995 9509
rect 23937 9469 23949 9503
rect 23983 9500 23995 9503
rect 24210 9500 24216 9512
rect 23983 9472 24216 9500
rect 23983 9469 23995 9472
rect 23937 9463 23995 9469
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9500 24915 9503
rect 25498 9500 25504 9512
rect 24903 9472 25504 9500
rect 24903 9469 24915 9472
rect 24857 9463 24915 9469
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 26694 9500 26700 9512
rect 26655 9472 26700 9500
rect 26694 9460 26700 9472
rect 26752 9460 26758 9512
rect 19886 9392 19892 9444
rect 19944 9432 19950 9444
rect 20349 9435 20407 9441
rect 20349 9432 20361 9435
rect 19944 9404 20361 9432
rect 19944 9392 19950 9404
rect 20349 9401 20361 9404
rect 20395 9401 20407 9435
rect 20349 9395 20407 9401
rect 20441 9435 20499 9441
rect 20441 9401 20453 9435
rect 20487 9432 20499 9435
rect 21008 9432 21036 9460
rect 25130 9441 25136 9444
rect 20487 9404 21036 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 25124 9395 25136 9441
rect 25188 9432 25194 9444
rect 25188 9404 25224 9432
rect 25130 9392 25136 9395
rect 25188 9392 25194 9404
rect 21542 9364 21548 9376
rect 19720 9336 21548 9364
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 23014 9324 23020 9376
rect 23072 9364 23078 9376
rect 23566 9364 23572 9376
rect 23072 9336 23572 9364
rect 23072 9324 23078 9336
rect 23566 9324 23572 9336
rect 23624 9324 23630 9376
rect 25038 9324 25044 9376
rect 25096 9364 25102 9376
rect 26237 9367 26295 9373
rect 26237 9364 26249 9367
rect 25096 9336 26249 9364
rect 25096 9324 25102 9336
rect 26237 9333 26249 9336
rect 26283 9333 26295 9367
rect 26237 9327 26295 9333
rect 1104 9274 28428 9296
rect 1104 9222 10090 9274
rect 10142 9222 10154 9274
rect 10206 9222 10218 9274
rect 10270 9222 10282 9274
rect 10334 9222 19198 9274
rect 19250 9222 19262 9274
rect 19314 9222 19326 9274
rect 19378 9222 19390 9274
rect 19442 9222 28428 9274
rect 1104 9200 28428 9222
rect 2682 9160 2688 9172
rect 2643 9132 2688 9160
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4890 9160 4896 9172
rect 4479 9132 4896 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5169 9163 5227 9169
rect 5169 9129 5181 9163
rect 5215 9160 5227 9163
rect 5258 9160 5264 9172
rect 5215 9132 5264 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 6914 9160 6920 9172
rect 6472 9132 6776 9160
rect 6875 9132 6920 9160
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2774 9092 2780 9104
rect 2455 9064 2780 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 2774 9052 2780 9064
rect 2832 9052 2838 9104
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 3660 9064 5120 9092
rect 3660 9052 3666 9064
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 2133 9027 2191 9033
rect 2133 9024 2145 9027
rect 2096 8996 2145 9024
rect 2096 8984 2102 8996
rect 2133 8993 2145 8996
rect 2179 8993 2191 9027
rect 2133 8987 2191 8993
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 8993 2375 9027
rect 2317 8987 2375 8993
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 8993 2559 9027
rect 2792 9024 2820 9052
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 2792 8996 3157 9024
rect 2501 8987 2559 8993
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 2332 8888 2360 8987
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 2516 8956 2544 8987
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 5092 9033 5120 9064
rect 5350 9052 5356 9104
rect 5408 9092 5414 9104
rect 5408 9064 6408 9092
rect 5408 9052 5414 9064
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 4304 8996 4353 9024
rect 4304 8984 4310 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 5994 9024 6000 9036
rect 5951 8996 6000 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6380 9033 6408 9064
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 8993 6423 9027
rect 6472 9024 6500 9132
rect 6638 9092 6644 9104
rect 6599 9064 6644 9092
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 6748 9092 6776 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7834 9160 7840 9172
rect 7432 9132 7840 9160
rect 7432 9120 7438 9132
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 9508 9132 9895 9160
rect 7208 9092 7236 9120
rect 7466 9092 7472 9104
rect 6748 9064 7472 9092
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 9122 9092 9128 9104
rect 8036 9064 9128 9092
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 6472 8996 6561 9024
rect 6365 8987 6423 8993
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 6730 9024 6736 9036
rect 6691 8996 6736 9024
rect 6549 8987 6607 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 8036 9033 8064 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7248 8996 7573 9024
rect 7248 8984 7254 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 9024 8447 9027
rect 9214 9024 9220 9036
rect 8435 8996 9220 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 9508 9033 9536 9132
rect 9628 9052 9634 9104
rect 9686 9101 9692 9104
rect 9686 9095 9735 9101
rect 9686 9061 9689 9095
rect 9723 9061 9735 9095
rect 9867 9092 9895 9132
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 10778 9160 10784 9172
rect 10468 9132 10784 9160
rect 10468 9120 10474 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 16761 9163 16819 9169
rect 16761 9160 16773 9163
rect 13780 9132 16773 9160
rect 13780 9120 13786 9132
rect 16761 9129 16773 9132
rect 16807 9129 16819 9163
rect 20530 9160 20536 9172
rect 20491 9132 20536 9160
rect 16761 9123 16819 9129
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 23256 9132 23305 9160
rect 23256 9120 23262 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 24210 9160 24216 9172
rect 24171 9132 24216 9160
rect 23293 9123 23351 9129
rect 24210 9120 24216 9132
rect 24268 9120 24274 9172
rect 25590 9120 25596 9172
rect 25648 9160 25654 9172
rect 25777 9163 25835 9169
rect 25777 9160 25789 9163
rect 25648 9132 25789 9160
rect 25648 9120 25654 9132
rect 25777 9129 25789 9132
rect 25823 9129 25835 9163
rect 25777 9123 25835 9129
rect 26418 9120 26424 9172
rect 26476 9160 26482 9172
rect 26973 9163 27031 9169
rect 26973 9160 26985 9163
rect 26476 9132 26985 9160
rect 26476 9120 26482 9132
rect 26973 9129 26985 9132
rect 27019 9129 27031 9163
rect 26973 9123 27031 9129
rect 10965 9095 11023 9101
rect 10965 9092 10977 9095
rect 9867 9064 10977 9092
rect 9686 9055 9735 9061
rect 10965 9061 10977 9064
rect 11011 9061 11023 9095
rect 12713 9095 12771 9101
rect 10965 9055 11023 9061
rect 11532 9064 12020 9092
rect 9686 9052 9692 9055
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9777 9027 9835 9033
rect 9777 8993 9789 9027
rect 9823 8993 9835 9027
rect 9777 8987 9835 8993
rect 9907 9027 9965 9033
rect 9907 8993 9919 9027
rect 9953 9024 9965 9027
rect 10042 9024 10048 9036
rect 9953 8996 10048 9024
rect 9953 8993 9965 8996
rect 9907 8987 9965 8993
rect 2464 8928 2544 8956
rect 3237 8959 3295 8965
rect 2464 8916 2470 8928
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 3283 8928 7757 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 7892 8928 8309 8956
rect 7892 8916 7898 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 9784 8956 9812 8987
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10870 9024 10876 9036
rect 10831 8996 10876 9024
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11054 9024 11060 9036
rect 11015 8996 11060 9024
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11330 9024 11336 9036
rect 11243 8996 11336 9024
rect 11330 8984 11336 8996
rect 11388 9024 11394 9036
rect 11532 9024 11560 9064
rect 11388 8996 11560 9024
rect 11388 8984 11394 8996
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11664 8996 11713 9024
rect 11664 8984 11670 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 11701 8987 11759 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 11992 9024 12020 9064
rect 12713 9061 12725 9095
rect 12759 9092 12771 9095
rect 15010 9092 15016 9104
rect 12759 9064 14872 9092
rect 14971 9064 15016 9092
rect 12759 9061 12771 9064
rect 12713 9055 12771 9061
rect 12894 9024 12900 9036
rect 11992 8996 12900 9024
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 9024 13415 9027
rect 13446 9024 13452 9036
rect 13403 8996 13452 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 10410 8956 10416 8968
rect 9784 8928 10416 8956
rect 8297 8919 8355 8925
rect 10410 8916 10416 8928
rect 10468 8956 10474 8968
rect 13630 8956 13636 8968
rect 10468 8928 13636 8956
rect 10468 8916 10474 8928
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 2332 8860 2774 8888
rect 2746 8820 2774 8860
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5350 8888 5356 8900
rect 5040 8860 5356 8888
rect 5040 8848 5046 8860
rect 5350 8848 5356 8860
rect 5408 8888 5414 8900
rect 5721 8891 5779 8897
rect 5721 8888 5733 8891
rect 5408 8860 5733 8888
rect 5408 8848 5414 8860
rect 5721 8857 5733 8860
rect 5767 8857 5779 8891
rect 5721 8851 5779 8857
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 14752 8888 14780 8987
rect 8251 8860 14780 8888
rect 14844 8888 14872 9064
rect 15010 9052 15016 9064
rect 15068 9052 15074 9104
rect 15654 9052 15660 9104
rect 15712 9092 15718 9104
rect 15712 9064 17080 9092
rect 15712 9052 15718 9064
rect 14918 8984 14924 9036
rect 14976 9024 14982 9036
rect 15105 9027 15163 9033
rect 14976 8996 15021 9024
rect 14976 8984 14982 8996
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 16298 9024 16304 9036
rect 15151 8996 16304 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 16574 9024 16580 9036
rect 16535 8996 16580 9024
rect 16574 8984 16580 8996
rect 16632 9024 16638 9036
rect 16942 9024 16948 9036
rect 16632 8996 16948 9024
rect 16632 8984 16638 8996
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17052 9024 17080 9064
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 17681 9095 17739 9101
rect 17681 9092 17693 9095
rect 17276 9064 17693 9092
rect 17276 9052 17282 9064
rect 17681 9061 17693 9064
rect 17727 9061 17739 9095
rect 17681 9055 17739 9061
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 19886 9092 19892 9104
rect 17828 9064 19892 9092
rect 17828 9052 17834 9064
rect 19886 9052 19892 9064
rect 19944 9092 19950 9104
rect 20165 9095 20223 9101
rect 20165 9092 20177 9095
rect 19944 9064 20177 9092
rect 19944 9052 19950 9064
rect 20165 9061 20177 9064
rect 20211 9061 20223 9095
rect 20165 9055 20223 9061
rect 20257 9095 20315 9101
rect 20257 9061 20269 9095
rect 20303 9092 20315 9095
rect 20438 9092 20444 9104
rect 20303 9064 20444 9092
rect 20303 9061 20315 9064
rect 20257 9055 20315 9061
rect 20438 9052 20444 9064
rect 20496 9052 20502 9104
rect 22094 9052 22100 9104
rect 22152 9092 22158 9104
rect 22925 9095 22983 9101
rect 22925 9092 22937 9095
rect 22152 9064 22937 9092
rect 22152 9052 22158 9064
rect 22925 9061 22937 9064
rect 22971 9092 22983 9095
rect 25409 9095 25467 9101
rect 25409 9092 25421 9095
rect 22971 9064 25421 9092
rect 22971 9061 22983 9064
rect 22925 9055 22983 9061
rect 25409 9061 25421 9064
rect 25455 9061 25467 9095
rect 25409 9055 25467 9061
rect 25501 9095 25559 9101
rect 25501 9061 25513 9095
rect 25547 9092 25559 9095
rect 26142 9092 26148 9104
rect 25547 9064 26148 9092
rect 25547 9061 25559 9064
rect 25501 9055 25559 9061
rect 18417 9027 18475 9033
rect 18417 9024 18429 9027
rect 17052 8996 18429 9024
rect 18417 8993 18429 8996
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 19794 8984 19800 9036
rect 19852 9024 19858 9036
rect 19981 9027 20039 9033
rect 19981 9024 19993 9027
rect 19852 8996 19993 9024
rect 19852 8984 19858 8996
rect 19981 8993 19993 8996
rect 20027 8993 20039 9027
rect 19981 8987 20039 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 15746 8916 15752 8968
rect 15804 8956 15810 8968
rect 19886 8956 19892 8968
rect 15804 8928 19892 8956
rect 15804 8916 15810 8928
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 17586 8888 17592 8900
rect 14844 8860 17592 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 17586 8848 17592 8860
rect 17644 8848 17650 8900
rect 17862 8888 17868 8900
rect 17823 8860 17868 8888
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 19702 8888 19708 8900
rect 17972 8860 19708 8888
rect 5902 8820 5908 8832
rect 2746 8792 5908 8820
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 10045 8823 10103 8829
rect 10045 8820 10057 8823
rect 8536 8792 10057 8820
rect 8536 8780 8542 8792
rect 10045 8789 10057 8792
rect 10091 8789 10103 8823
rect 10045 8783 10103 8789
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11606 8820 11612 8832
rect 10836 8792 11612 8820
rect 10836 8780 10842 8792
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 12952 8792 13553 8820
rect 12952 8780 12958 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 13541 8783 13599 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 17770 8820 17776 8832
rect 16908 8792 17776 8820
rect 16908 8780 16914 8792
rect 17770 8780 17776 8792
rect 17828 8820 17834 8832
rect 17972 8820 18000 8860
rect 19702 8848 19708 8860
rect 19760 8848 19766 8900
rect 19996 8888 20024 8987
rect 20364 8956 20392 8987
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 22741 9027 22799 9033
rect 22741 9024 22753 9027
rect 21876 8996 22753 9024
rect 21876 8984 21882 8996
rect 22741 8993 22753 8996
rect 22787 8993 22799 9027
rect 23014 9024 23020 9036
rect 22975 8996 23020 9024
rect 22741 8987 22799 8993
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 23109 9027 23167 9033
rect 23109 8993 23121 9027
rect 23155 8993 23167 9027
rect 23109 8987 23167 8993
rect 24121 9027 24179 9033
rect 24121 8993 24133 9027
rect 24167 9024 24179 9027
rect 25038 9024 25044 9036
rect 24167 8996 25044 9024
rect 24167 8993 24179 8996
rect 24121 8987 24179 8993
rect 21910 8956 21916 8968
rect 20364 8928 21916 8956
rect 21910 8916 21916 8928
rect 21968 8956 21974 8968
rect 23124 8956 23152 8987
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 25225 9027 25283 9033
rect 25225 8993 25237 9027
rect 25271 9024 25283 9027
rect 25314 9024 25320 9036
rect 25271 8996 25320 9024
rect 25271 8993 25283 8996
rect 25225 8987 25283 8993
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 25424 8968 25452 9055
rect 26142 9052 26148 9064
rect 26200 9052 26206 9104
rect 25617 9027 25675 9033
rect 25617 9024 25629 9027
rect 25608 8993 25629 9024
rect 25663 8993 25675 9027
rect 26786 9024 26792 9036
rect 26747 8996 26792 9024
rect 25608 8987 25675 8993
rect 21968 8928 23152 8956
rect 21968 8916 21974 8928
rect 25406 8916 25412 8968
rect 25464 8916 25470 8968
rect 21818 8888 21824 8900
rect 19996 8860 21824 8888
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 25608 8888 25636 8987
rect 26786 8984 26792 8996
rect 26844 8984 26850 9036
rect 27522 9024 27528 9036
rect 27483 8996 27528 9024
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 27706 8888 27712 8900
rect 24964 8860 25636 8888
rect 27667 8860 27712 8888
rect 24964 8832 24992 8860
rect 27706 8848 27712 8860
rect 27764 8848 27770 8900
rect 18506 8820 18512 8832
rect 17828 8792 18000 8820
rect 18467 8792 18512 8820
rect 17828 8780 17834 8792
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 18690 8780 18696 8832
rect 18748 8820 18754 8832
rect 19610 8820 19616 8832
rect 18748 8792 19616 8820
rect 18748 8780 18754 8792
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 22002 8780 22008 8832
rect 22060 8820 22066 8832
rect 24946 8820 24952 8832
rect 22060 8792 24952 8820
rect 22060 8780 22066 8792
rect 24946 8780 24952 8792
rect 25004 8780 25010 8832
rect 1104 8730 28428 8752
rect 1104 8678 5536 8730
rect 5588 8678 5600 8730
rect 5652 8678 5664 8730
rect 5716 8678 5728 8730
rect 5780 8678 14644 8730
rect 14696 8678 14708 8730
rect 14760 8678 14772 8730
rect 14824 8678 14836 8730
rect 14888 8678 23752 8730
rect 23804 8678 23816 8730
rect 23868 8678 23880 8730
rect 23932 8678 23944 8730
rect 23996 8678 28428 8730
rect 1104 8656 28428 8678
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 4065 8619 4123 8625
rect 4065 8585 4077 8619
rect 4111 8616 4123 8619
rect 4154 8616 4160 8628
rect 4111 8588 4160 8616
rect 4111 8585 4123 8588
rect 4065 8579 4123 8585
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 4706 8616 4712 8628
rect 4387 8588 4712 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 7653 8619 7711 8625
rect 7653 8585 7665 8619
rect 7699 8616 7711 8619
rect 7834 8616 7840 8628
rect 7699 8588 7840 8616
rect 7699 8585 7711 8588
rect 7653 8579 7711 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 8220 8588 9597 8616
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 8220 8548 8248 8588
rect 9585 8585 9597 8588
rect 9631 8616 9643 8619
rect 10042 8616 10048 8628
rect 9631 8588 10048 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 11330 8616 11336 8628
rect 10520 8588 11336 8616
rect 5224 8520 8248 8548
rect 5224 8508 5230 8520
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 10520 8548 10548 8588
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 15746 8616 15752 8628
rect 13740 8588 15752 8616
rect 9272 8520 10548 8548
rect 9272 8508 9278 8520
rect 2406 8440 2412 8492
rect 2464 8480 2470 8492
rect 2464 8452 2728 8480
rect 2464 8440 2470 8452
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 2096 8384 2329 8412
rect 2096 8372 2102 8384
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2498 8412 2504 8424
rect 2459 8384 2504 8412
rect 2317 8375 2375 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2700 8421 2728 8452
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 9456 8452 10241 8480
rect 9456 8440 9462 8452
rect 10229 8449 10241 8452
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8381 2743 8415
rect 3878 8412 3884 8424
rect 3839 8384 3884 8412
rect 2685 8375 2743 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8294 8412 8300 8424
rect 8251 8384 8300 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8478 8421 8484 8424
rect 8472 8412 8484 8421
rect 8439 8384 8484 8412
rect 8472 8375 8484 8384
rect 8478 8372 8484 8375
rect 8536 8372 8542 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10520 8421 10548 8520
rect 10781 8551 10839 8557
rect 10781 8517 10793 8551
rect 10827 8517 10839 8551
rect 10781 8511 10839 8517
rect 10796 8480 10824 8511
rect 10796 8452 13400 8480
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 9732 8384 10057 8412
rect 9732 8372 9738 8384
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10045 8375 10103 8381
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 10836 8384 10885 8412
rect 10836 8372 10842 8384
rect 10873 8381 10885 8384
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8381 11023 8415
rect 12066 8412 12072 8424
rect 12027 8384 12072 8412
rect 10965 8375 11023 8381
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 3602 8344 3608 8356
rect 2639 8316 3608 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 3602 8304 3608 8316
rect 3660 8304 3666 8356
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 10980 8344 11008 8375
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 12216 8384 12357 8412
rect 12216 8372 12222 8384
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12526 8412 12532 8424
rect 12483 8384 12532 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 13372 8421 13400 8452
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13630 8412 13636 8424
rect 13591 8384 13636 8412
rect 13357 8375 13415 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13740 8421 13768 8588
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18966 8616 18972 8628
rect 18279 8588 18972 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 20162 8616 20168 8628
rect 20123 8588 20168 8616
rect 20162 8576 20168 8588
rect 20220 8576 20226 8628
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 23198 8616 23204 8628
rect 22796 8588 23204 8616
rect 22796 8576 22802 8588
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 25130 8616 25136 8628
rect 25091 8588 25136 8616
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 17589 8551 17647 8557
rect 17589 8517 17601 8551
rect 17635 8548 17647 8551
rect 17770 8548 17776 8560
rect 17635 8520 17776 8548
rect 17635 8517 17647 8520
rect 17589 8511 17647 8517
rect 13924 8480 13952 8511
rect 17770 8508 17776 8520
rect 17828 8508 17834 8560
rect 20254 8508 20260 8560
rect 20312 8548 20318 8560
rect 25314 8548 25320 8560
rect 20312 8520 25320 8548
rect 20312 8508 20318 8520
rect 13924 8452 14504 8480
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 14366 8412 14372 8424
rect 14327 8384 14372 8412
rect 13725 8375 13783 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14476 8412 14504 8452
rect 20070 8440 20076 8492
rect 20128 8480 20134 8492
rect 20128 8452 21588 8480
rect 20128 8440 20134 8452
rect 14625 8415 14683 8421
rect 14625 8412 14637 8415
rect 14476 8384 14637 8412
rect 14625 8381 14637 8384
rect 14671 8381 14683 8415
rect 14625 8375 14683 8381
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 17218 8412 17224 8424
rect 15620 8384 17224 8412
rect 15620 8372 15626 8384
rect 17218 8372 17224 8384
rect 17276 8412 17282 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 17276 8384 17417 8412
rect 17276 8372 17282 8384
rect 17405 8381 17417 8384
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 18046 8372 18052 8424
rect 18104 8412 18110 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 18104 8384 18153 8412
rect 18104 8372 18110 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 19058 8421 19064 8424
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18748 8384 18797 8412
rect 18748 8372 18754 8384
rect 18785 8381 18797 8384
rect 18831 8381 18843 8415
rect 18785 8375 18843 8381
rect 19052 8375 19064 8421
rect 19116 8412 19122 8424
rect 19116 8384 19152 8412
rect 19058 8372 19064 8375
rect 19116 8372 19122 8384
rect 20162 8372 20168 8424
rect 20220 8412 20226 8424
rect 21560 8421 21588 8452
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20220 8384 20729 8412
rect 20220 8372 20226 8384
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 21545 8415 21603 8421
rect 21545 8381 21557 8415
rect 21591 8381 21603 8415
rect 21545 8375 21603 8381
rect 21726 8372 21732 8424
rect 21784 8412 21790 8424
rect 22741 8415 22799 8421
rect 22741 8412 22753 8415
rect 21784 8384 22753 8412
rect 21784 8372 21790 8384
rect 22741 8381 22753 8384
rect 22787 8412 22799 8415
rect 23474 8412 23480 8424
rect 22787 8384 23480 8412
rect 22787 8381 22799 8384
rect 22741 8375 22799 8381
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8412 24179 8415
rect 24394 8412 24400 8424
rect 24167 8384 24400 8412
rect 24167 8381 24179 8384
rect 24121 8375 24179 8381
rect 24394 8372 24400 8384
rect 24452 8372 24458 8424
rect 24596 8421 24624 8520
rect 25314 8508 25320 8520
rect 25372 8508 25378 8560
rect 26145 8551 26203 8557
rect 26145 8517 26157 8551
rect 26191 8548 26203 8551
rect 26234 8548 26240 8560
rect 26191 8520 26240 8548
rect 26191 8517 26203 8520
rect 26145 8511 26203 8517
rect 26234 8508 26240 8520
rect 26292 8508 26298 8560
rect 25038 8480 25044 8492
rect 24872 8452 25044 8480
rect 24872 8421 24900 8452
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 24581 8415 24639 8421
rect 24581 8381 24593 8415
rect 24627 8381 24639 8415
rect 24581 8375 24639 8381
rect 24857 8415 24915 8421
rect 24857 8381 24869 8415
rect 24903 8381 24915 8415
rect 24857 8375 24915 8381
rect 24946 8372 24952 8424
rect 25004 8412 25010 8424
rect 25004 8384 25049 8412
rect 25004 8372 25010 8384
rect 25130 8372 25136 8424
rect 25188 8412 25194 8424
rect 25593 8415 25651 8421
rect 25593 8412 25605 8415
rect 25188 8384 25605 8412
rect 25188 8372 25194 8384
rect 25593 8381 25605 8384
rect 25639 8381 25651 8415
rect 25866 8412 25872 8424
rect 25827 8384 25872 8412
rect 25593 8375 25651 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 25961 8415 26019 8421
rect 25961 8381 25973 8415
rect 26007 8381 26019 8415
rect 26694 8412 26700 8424
rect 26655 8384 26700 8412
rect 25961 8375 26019 8381
rect 8812 8316 11008 8344
rect 8812 8304 8818 8316
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11974 8344 11980 8356
rect 11112 8316 11980 8344
rect 11112 8304 11118 8316
rect 11974 8304 11980 8316
rect 12032 8344 12038 8356
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 12032 8316 12265 8344
rect 12032 8304 12038 8316
rect 12253 8313 12265 8316
rect 12299 8313 12311 8347
rect 13538 8344 13544 8356
rect 13499 8316 13544 8344
rect 12253 8307 12311 8313
rect 13538 8304 13544 8316
rect 13596 8344 13602 8356
rect 14182 8344 14188 8356
rect 13596 8316 14188 8344
rect 13596 8304 13602 8316
rect 14182 8304 14188 8316
rect 14240 8304 14246 8356
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 17644 8316 21404 8344
rect 17644 8304 17650 8316
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7006 8276 7012 8288
rect 6963 8248 7012 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 12618 8276 12624 8288
rect 12579 8248 12624 8276
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 20714 8276 20720 8288
rect 18748 8248 20720 8276
rect 18748 8236 18754 8248
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 20809 8279 20867 8285
rect 20809 8245 20821 8279
rect 20855 8276 20867 8279
rect 21174 8276 21180 8288
rect 20855 8248 21180 8276
rect 20855 8245 20867 8248
rect 20809 8239 20867 8245
rect 21174 8236 21180 8248
rect 21232 8236 21238 8288
rect 21376 8285 21404 8316
rect 22186 8304 22192 8356
rect 22244 8344 22250 8356
rect 24765 8347 24823 8353
rect 24765 8344 24777 8347
rect 22244 8316 24777 8344
rect 22244 8304 22250 8316
rect 24765 8313 24777 8316
rect 24811 8344 24823 8347
rect 25777 8347 25835 8353
rect 25777 8344 25789 8347
rect 24811 8316 25789 8344
rect 24811 8313 24823 8316
rect 24765 8307 24823 8313
rect 25777 8313 25789 8316
rect 25823 8313 25835 8347
rect 25777 8307 25835 8313
rect 21361 8279 21419 8285
rect 21361 8245 21373 8279
rect 21407 8245 21419 8279
rect 21361 8239 21419 8245
rect 22833 8279 22891 8285
rect 22833 8245 22845 8279
rect 22879 8276 22891 8279
rect 23106 8276 23112 8288
rect 22879 8248 23112 8276
rect 22879 8245 22891 8248
rect 22833 8239 22891 8245
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 23937 8279 23995 8285
rect 23937 8245 23949 8279
rect 23983 8276 23995 8279
rect 24946 8276 24952 8288
rect 23983 8248 24952 8276
rect 23983 8245 23995 8248
rect 23937 8239 23995 8245
rect 24946 8236 24952 8248
rect 25004 8276 25010 8288
rect 25498 8276 25504 8288
rect 25004 8248 25504 8276
rect 25004 8236 25010 8248
rect 25498 8236 25504 8248
rect 25556 8236 25562 8288
rect 25590 8236 25596 8288
rect 25648 8276 25654 8288
rect 25976 8276 26004 8375
rect 26694 8372 26700 8384
rect 26752 8372 26758 8424
rect 26878 8276 26884 8288
rect 25648 8248 26004 8276
rect 26839 8248 26884 8276
rect 25648 8236 25654 8248
rect 26878 8236 26884 8248
rect 26936 8236 26942 8288
rect 1104 8186 28428 8208
rect 1104 8134 10090 8186
rect 10142 8134 10154 8186
rect 10206 8134 10218 8186
rect 10270 8134 10282 8186
rect 10334 8134 19198 8186
rect 19250 8134 19262 8186
rect 19314 8134 19326 8186
rect 19378 8134 19390 8186
rect 19442 8134 28428 8186
rect 1104 8112 28428 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1544 8044 1593 8072
rect 1544 8032 1550 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 1581 8035 1639 8041
rect 6012 8044 7849 8072
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 5712 8007 5770 8013
rect 4755 7976 5672 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 1578 7896 1584 7948
rect 1636 7936 1642 7948
rect 2133 7939 2191 7945
rect 2133 7936 2145 7939
rect 1636 7908 2145 7936
rect 1636 7896 1642 7908
rect 2133 7905 2145 7908
rect 2179 7905 2191 7939
rect 4430 7936 4436 7948
rect 4391 7908 4436 7936
rect 2133 7899 2191 7905
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7905 4675 7939
rect 4617 7899 4675 7905
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 5074 7936 5080 7948
rect 4847 7908 5080 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 4632 7868 4660 7899
rect 5074 7896 5080 7908
rect 5132 7936 5138 7948
rect 5132 7908 5396 7936
rect 5132 7896 5138 7908
rect 5166 7868 5172 7880
rect 4632 7840 5172 7868
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 4982 7732 4988 7744
rect 4943 7704 4988 7732
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5368 7732 5396 7908
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5644 7936 5672 7976
rect 5712 7973 5724 8007
rect 5758 8004 5770 8007
rect 6012 8004 6040 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 8352 8044 9873 8072
rect 8352 8032 8358 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 5758 7976 6040 8004
rect 9876 8004 9904 8035
rect 12158 8032 12164 8084
rect 12216 8072 12222 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 12216 8044 13737 8072
rect 12216 8032 12222 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 15528 8044 17049 8072
rect 15528 8032 15534 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 18506 8072 18512 8084
rect 17037 8035 17095 8041
rect 17604 8044 18512 8072
rect 12618 8013 12624 8016
rect 12612 8004 12624 8013
rect 9876 7976 12388 8004
rect 12579 7976 12624 8004
rect 5758 7973 5770 7976
rect 5712 7967 5770 7973
rect 5994 7936 6000 7948
rect 5500 7908 5545 7936
rect 5644 7908 6000 7936
rect 5500 7896 5506 7908
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 6144 7908 7297 7936
rect 6144 7896 6150 7908
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 7466 7936 7472 7948
rect 7427 7908 7472 7936
rect 7285 7899 7343 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 7699 7908 7972 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 7576 7868 7604 7899
rect 7834 7868 7840 7880
rect 6840 7840 7840 7868
rect 6840 7809 6868 7840
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7769 6883 7803
rect 6825 7763 6883 7769
rect 7944 7732 7972 7908
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10520 7945 10548 7976
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 10008 7908 10057 7936
rect 10008 7896 10014 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10772 7939 10830 7945
rect 10772 7905 10784 7939
rect 10818 7936 10830 7939
rect 11330 7936 11336 7948
rect 10818 7908 11336 7936
rect 10818 7905 10830 7908
rect 10772 7899 10830 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 12360 7945 12388 7976
rect 12612 7967 12624 7976
rect 12618 7964 12624 7967
rect 12676 7964 12682 8016
rect 15004 8007 15062 8013
rect 15004 7973 15016 8007
rect 15050 8004 15062 8007
rect 15286 8004 15292 8016
rect 15050 7976 15292 8004
rect 15050 7973 15062 7976
rect 15004 7967 15062 7973
rect 15286 7964 15292 7976
rect 15344 7964 15350 8016
rect 17604 8004 17632 8044
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 20349 8075 20407 8081
rect 20349 8072 20361 8075
rect 19024 8044 20361 8072
rect 19024 8032 19030 8044
rect 20349 8041 20361 8044
rect 20395 8041 20407 8075
rect 20349 8035 20407 8041
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21177 8075 21235 8081
rect 21177 8072 21189 8075
rect 21140 8044 21189 8072
rect 21140 8032 21146 8044
rect 21177 8041 21189 8044
rect 21223 8041 21235 8075
rect 21177 8035 21235 8041
rect 22922 8032 22928 8084
rect 22980 8072 22986 8084
rect 23385 8075 23443 8081
rect 23385 8072 23397 8075
rect 22980 8044 23397 8072
rect 22980 8032 22986 8044
rect 23385 8041 23397 8044
rect 23431 8041 23443 8075
rect 25774 8072 25780 8084
rect 23385 8035 23443 8041
rect 23952 8044 25780 8072
rect 21729 8007 21787 8013
rect 21729 8004 21741 8007
rect 17512 7976 17632 8004
rect 17880 7976 18920 8004
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 13078 7936 13084 7948
rect 12391 7908 13084 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 13078 7896 13084 7908
rect 13136 7936 13142 7948
rect 14366 7936 14372 7948
rect 13136 7908 14372 7936
rect 13136 7896 13142 7908
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 14424 7908 14749 7936
rect 14424 7896 14430 7908
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 16574 7936 16580 7948
rect 16535 7908 16580 7936
rect 14737 7899 14795 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 17512 7945 17540 7976
rect 17880 7948 17908 7976
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17678 7936 17684 7948
rect 17591 7908 17684 7936
rect 17497 7899 17555 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17696 7868 17724 7896
rect 17184 7840 17724 7868
rect 17788 7868 17816 7899
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 18506 7936 18512 7948
rect 17920 7908 17965 7936
rect 18467 7908 18512 7936
rect 17920 7896 17926 7908
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 18690 7936 18696 7948
rect 18651 7908 18696 7936
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 18892 7945 18920 7976
rect 20548 7976 21741 8004
rect 18785 7939 18843 7945
rect 18785 7905 18797 7939
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 18966 7936 18972 7948
rect 18923 7908 18972 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 18046 7868 18052 7880
rect 17788 7840 18052 7868
rect 17184 7828 17190 7840
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18800 7868 18828 7899
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 20070 7896 20076 7948
rect 20128 7936 20134 7948
rect 20441 7939 20499 7945
rect 20441 7936 20453 7939
rect 20128 7908 20453 7936
rect 20128 7896 20134 7908
rect 20441 7905 20453 7908
rect 20487 7905 20499 7939
rect 20548 7936 20576 7976
rect 21729 7973 21741 7976
rect 21775 7973 21787 8007
rect 21729 7967 21787 7973
rect 21818 7964 21824 8016
rect 21876 8004 21882 8016
rect 23952 8004 23980 8044
rect 25774 8032 25780 8044
rect 25832 8032 25838 8084
rect 25958 8032 25964 8084
rect 26016 8072 26022 8084
rect 27341 8075 27399 8081
rect 27341 8072 27353 8075
rect 26016 8044 27353 8072
rect 26016 8032 26022 8044
rect 27341 8041 27353 8044
rect 27387 8041 27399 8075
rect 27341 8035 27399 8041
rect 25976 8004 26004 8032
rect 26234 8013 26240 8016
rect 26228 8004 26240 8013
rect 21876 7976 23980 8004
rect 24136 7976 26004 8004
rect 26195 7976 26240 8004
rect 21876 7964 21882 7976
rect 20898 7945 20904 7948
rect 20625 7939 20683 7945
rect 20625 7936 20637 7939
rect 20548 7908 20637 7936
rect 20441 7899 20499 7905
rect 20625 7905 20637 7908
rect 20671 7905 20683 7939
rect 20855 7939 20904 7945
rect 20855 7936 20867 7939
rect 20811 7908 20867 7936
rect 20625 7899 20683 7905
rect 20855 7905 20867 7908
rect 20901 7905 20904 7939
rect 20855 7899 20904 7905
rect 20898 7896 20904 7899
rect 20956 7896 20962 7948
rect 20993 7939 21051 7945
rect 20993 7905 21005 7939
rect 21039 7936 21051 7939
rect 21174 7936 21180 7948
rect 21039 7908 21180 7936
rect 21039 7905 21051 7908
rect 20993 7899 21051 7905
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 21637 7939 21695 7945
rect 21637 7905 21649 7939
rect 21683 7936 21695 7939
rect 22094 7936 22100 7948
rect 21683 7908 22100 7936
rect 21683 7905 21695 7908
rect 21637 7899 21695 7905
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7905 22707 7939
rect 22830 7936 22836 7948
rect 22791 7908 22836 7936
rect 22649 7899 22707 7905
rect 20162 7868 20168 7880
rect 18800 7840 20168 7868
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20717 7871 20775 7877
rect 20717 7868 20729 7871
rect 20395 7840 20729 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20717 7837 20729 7840
rect 20763 7837 20775 7871
rect 20907 7868 20935 7896
rect 20717 7831 20775 7837
rect 20824 7840 20935 7868
rect 16390 7760 16396 7812
rect 16448 7800 16454 7812
rect 20824 7800 20852 7840
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 22664 7868 22692 7899
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 23014 7936 23020 7948
rect 22975 7908 23020 7936
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 24136 7945 24164 7976
rect 26228 7967 26240 7976
rect 26234 7964 26240 7967
rect 26292 7964 26298 8016
rect 23201 7939 23259 7945
rect 23201 7905 23213 7939
rect 23247 7905 23259 7939
rect 23201 7899 23259 7905
rect 24121 7939 24179 7945
rect 24121 7905 24133 7939
rect 24167 7905 24179 7939
rect 24121 7899 24179 7905
rect 22738 7868 22744 7880
rect 21324 7840 22416 7868
rect 22664 7840 22744 7868
rect 21324 7828 21330 7840
rect 16448 7772 20852 7800
rect 22388 7800 22416 7840
rect 22738 7828 22744 7840
rect 22796 7828 22802 7880
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7837 22983 7871
rect 23216 7868 23244 7899
rect 24854 7896 24860 7948
rect 24912 7936 24918 7948
rect 25225 7939 25283 7945
rect 25225 7936 25237 7939
rect 24912 7908 25237 7936
rect 24912 7896 24918 7908
rect 25225 7905 25237 7908
rect 25271 7936 25283 7939
rect 25498 7936 25504 7948
rect 25271 7908 25504 7936
rect 25271 7905 25283 7908
rect 25225 7899 25283 7905
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 24213 7871 24271 7877
rect 24213 7868 24225 7871
rect 23216 7840 24225 7868
rect 22925 7831 22983 7837
rect 24213 7837 24225 7840
rect 24259 7837 24271 7871
rect 24213 7831 24271 7837
rect 22943 7800 22971 7831
rect 24946 7828 24952 7880
rect 25004 7868 25010 7880
rect 25961 7871 26019 7877
rect 25961 7868 25973 7871
rect 25004 7840 25973 7868
rect 25004 7828 25010 7840
rect 25961 7837 25973 7840
rect 26007 7837 26019 7871
rect 25961 7831 26019 7837
rect 22388 7772 22971 7800
rect 16448 7760 16454 7772
rect 5368 7704 7972 7732
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 11885 7735 11943 7741
rect 11885 7732 11897 7735
rect 11204 7704 11897 7732
rect 11204 7692 11210 7704
rect 11885 7701 11897 7704
rect 11931 7732 11943 7735
rect 12250 7732 12256 7744
rect 11931 7704 12256 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 16117 7735 16175 7741
rect 16117 7701 16129 7735
rect 16163 7732 16175 7735
rect 16298 7732 16304 7744
rect 16163 7704 16304 7732
rect 16163 7701 16175 7704
rect 16117 7695 16175 7701
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16853 7735 16911 7741
rect 16853 7701 16865 7735
rect 16899 7732 16911 7735
rect 17770 7732 17776 7744
rect 16899 7704 17776 7732
rect 16899 7701 16911 7704
rect 16853 7695 16911 7701
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 18012 7704 18061 7732
rect 18012 7692 18018 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 19058 7732 19064 7744
rect 19019 7704 19064 7732
rect 18049 7695 18107 7701
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 20349 7735 20407 7741
rect 20349 7701 20361 7735
rect 20395 7732 20407 7735
rect 22830 7732 22836 7744
rect 20395 7704 22836 7732
rect 20395 7701 20407 7704
rect 20349 7695 20407 7701
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 24210 7692 24216 7744
rect 24268 7732 24274 7744
rect 24762 7732 24768 7744
rect 24268 7704 24768 7732
rect 24268 7692 24274 7704
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 25314 7732 25320 7744
rect 25275 7704 25320 7732
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 1104 7642 28428 7664
rect 1104 7590 5536 7642
rect 5588 7590 5600 7642
rect 5652 7590 5664 7642
rect 5716 7590 5728 7642
rect 5780 7590 14644 7642
rect 14696 7590 14708 7642
rect 14760 7590 14772 7642
rect 14824 7590 14836 7642
rect 14888 7590 23752 7642
rect 23804 7590 23816 7642
rect 23868 7590 23880 7642
rect 23932 7590 23944 7642
rect 23996 7590 28428 7642
rect 1104 7568 28428 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 4062 7528 4068 7540
rect 3835 7500 4068 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 5350 7528 5356 7540
rect 4448 7500 5356 7528
rect 3970 7460 3976 7472
rect 3931 7432 3976 7460
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 2406 7392 2412 7404
rect 2148 7364 2412 7392
rect 1486 7324 1492 7336
rect 1447 7296 1492 7324
rect 1486 7284 1492 7296
rect 1544 7284 1550 7336
rect 2148 7333 2176 7364
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4448 7401 4476 7500
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 5994 7528 6000 7540
rect 5859 7500 6000 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 5994 7488 6000 7500
rect 6052 7528 6058 7540
rect 6822 7528 6828 7540
rect 6052 7500 6828 7528
rect 6052 7488 6058 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 10597 7531 10655 7537
rect 10597 7497 10609 7531
rect 10643 7528 10655 7531
rect 10870 7528 10876 7540
rect 10643 7500 10876 7528
rect 10643 7497 10655 7500
rect 10597 7491 10655 7497
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11940 7500 12173 7528
rect 11940 7488 11946 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 17034 7528 17040 7540
rect 16347 7500 17040 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17310 7488 17316 7540
rect 17368 7528 17374 7540
rect 19702 7528 19708 7540
rect 17368 7500 18736 7528
rect 19663 7500 19708 7528
rect 17368 7488 17374 7500
rect 7285 7463 7343 7469
rect 7285 7429 7297 7463
rect 7331 7460 7343 7463
rect 8110 7460 8116 7472
rect 7331 7432 8116 7460
rect 7331 7429 7343 7432
rect 7285 7423 7343 7429
rect 8110 7420 8116 7432
rect 8168 7460 8174 7472
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 8168 7432 11069 7460
rect 8168 7420 8174 7432
rect 11057 7429 11069 7432
rect 11103 7460 11115 7463
rect 12802 7460 12808 7472
rect 11103 7432 12808 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 12802 7420 12808 7432
rect 12860 7460 12866 7472
rect 13262 7460 13268 7472
rect 12860 7432 13268 7460
rect 12860 7420 12866 7432
rect 13262 7420 13268 7432
rect 13320 7420 13326 7472
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4212 7364 4445 7392
rect 4212 7352 4218 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7190 7392 7196 7404
rect 6871 7364 7196 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7650 7392 7656 7404
rect 7300 7364 7656 7392
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7293 2191 7327
rect 2314 7324 2320 7336
rect 2275 7296 2320 7324
rect 2133 7287 2191 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7324 2559 7327
rect 2866 7324 2872 7336
rect 2547 7296 2872 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 2866 7284 2872 7296
rect 2924 7324 2930 7336
rect 3535 7327 3593 7333
rect 2924 7296 3464 7324
rect 2924 7284 2930 7296
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 3142 7256 3148 7268
rect 2455 7228 3148 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 3436 7188 3464 7296
rect 3535 7293 3547 7327
rect 3581 7324 3593 7327
rect 4062 7324 4068 7336
rect 3581 7296 4068 7324
rect 3581 7293 3593 7296
rect 3535 7287 3593 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 4700 7327 4758 7333
rect 4700 7293 4712 7327
rect 4746 7324 4758 7327
rect 4982 7324 4988 7336
rect 4746 7296 4988 7324
rect 4746 7293 4758 7296
rect 4700 7287 4758 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5920 7324 5948 7352
rect 6546 7324 6552 7336
rect 5224 7296 6552 7324
rect 5224 7284 5230 7296
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 7006 7324 7012 7336
rect 6967 7296 7012 7324
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7300 7324 7328 7364
rect 7650 7352 7656 7364
rect 7708 7392 7714 7404
rect 8386 7392 8392 7404
rect 7708 7364 8392 7392
rect 7708 7352 7714 7364
rect 8386 7352 8392 7364
rect 8444 7392 8450 7404
rect 13354 7392 13360 7404
rect 8444 7364 10916 7392
rect 8444 7352 8450 7364
rect 7147 7296 7328 7324
rect 7377 7327 7435 7333
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7377 7293 7389 7327
rect 7423 7293 7435 7327
rect 7834 7324 7840 7336
rect 7795 7296 7840 7324
rect 7377 7287 7435 7293
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 7392 7256 7420 7287
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 10888 7333 10916 7364
rect 11164 7364 13360 7392
rect 11164 7333 11192 7364
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 17586 7352 17592 7404
rect 17644 7392 17650 7404
rect 17681 7395 17739 7401
rect 17681 7392 17693 7395
rect 17644 7364 17693 7392
rect 17644 7352 17650 7364
rect 17681 7361 17693 7364
rect 17727 7361 17739 7395
rect 18708 7392 18736 7500
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 20070 7528 20076 7540
rect 20031 7500 20076 7528
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 23293 7531 23351 7537
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 23382 7528 23388 7540
rect 23339 7500 23388 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 26237 7531 26295 7537
rect 26237 7528 26249 7531
rect 23532 7500 26249 7528
rect 23532 7488 23538 7500
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 19024 7432 21956 7460
rect 19024 7420 19030 7432
rect 21174 7392 21180 7404
rect 18708 7364 21180 7392
rect 17681 7355 17739 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 21818 7392 21824 7404
rect 21284 7364 21824 7392
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7324 12127 7327
rect 12158 7324 12164 7336
rect 12115 7296 12164 7324
rect 12115 7293 12127 7296
rect 12069 7287 12127 7293
rect 5960 7228 7420 7256
rect 10796 7256 10824 7287
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12308 7296 12725 7324
rect 12308 7284 12314 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 16482 7324 16488 7336
rect 16255 7296 16488 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 17954 7333 17960 7336
rect 17948 7324 17960 7333
rect 17915 7296 17960 7324
rect 17948 7287 17960 7296
rect 17954 7284 17960 7287
rect 18012 7284 18018 7336
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 19978 7324 19984 7336
rect 19659 7296 19984 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20530 7284 20536 7336
rect 20588 7324 20594 7336
rect 21284 7333 21312 7364
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 21928 7392 21956 7432
rect 22066 7432 23704 7460
rect 22066 7392 22094 7432
rect 22830 7392 22836 7404
rect 21928 7364 22094 7392
rect 22791 7364 22836 7392
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 23014 7392 23020 7404
rect 22971 7364 23020 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 23014 7352 23020 7364
rect 23072 7392 23078 7404
rect 23474 7392 23480 7404
rect 23072 7364 23480 7392
rect 23072 7352 23078 7364
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20588 7296 21097 7324
rect 20588 7284 20594 7296
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7293 21327 7327
rect 21450 7324 21456 7336
rect 21411 7296 21456 7324
rect 21269 7287 21327 7293
rect 21450 7284 21456 7296
rect 21508 7284 21514 7336
rect 22554 7324 22560 7336
rect 22515 7296 22560 7324
rect 22554 7284 22560 7296
rect 22612 7284 22618 7336
rect 22646 7284 22652 7336
rect 22704 7324 22710 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22704 7296 22753 7324
rect 22704 7284 22710 7296
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 23106 7324 23112 7336
rect 23067 7296 23112 7324
rect 22741 7287 22799 7293
rect 23106 7284 23112 7296
rect 23164 7284 23170 7336
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 10796 7228 12817 7256
rect 5960 7216 5966 7228
rect 12805 7225 12817 7228
rect 12851 7225 12863 7259
rect 12805 7219 12863 7225
rect 21361 7259 21419 7265
rect 21361 7225 21373 7259
rect 21407 7256 21419 7259
rect 22094 7256 22100 7268
rect 21407 7228 22100 7256
rect 21407 7225 21419 7228
rect 21361 7219 21419 7225
rect 22094 7216 22100 7228
rect 22152 7256 22158 7268
rect 22830 7256 22836 7268
rect 22152 7228 22836 7256
rect 22152 7216 22158 7228
rect 22830 7216 22836 7228
rect 22888 7216 22894 7268
rect 4706 7188 4712 7200
rect 3436 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 7929 7191 7987 7197
rect 7929 7188 7941 7191
rect 7432 7160 7941 7188
rect 7432 7148 7438 7160
rect 7929 7157 7941 7160
rect 7975 7157 7987 7191
rect 7929 7151 7987 7157
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 18046 7188 18052 7200
rect 8076 7160 18052 7188
rect 8076 7148 8082 7160
rect 18046 7148 18052 7160
rect 18104 7188 18110 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18104 7160 19073 7188
rect 18104 7148 18110 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 21637 7191 21695 7197
rect 21637 7157 21649 7191
rect 21683 7188 21695 7191
rect 22462 7188 22468 7200
rect 21683 7160 22468 7188
rect 21683 7157 21695 7160
rect 21637 7151 21695 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 23676 7188 23704 7432
rect 23842 7324 23848 7336
rect 23803 7296 23848 7324
rect 23842 7284 23848 7296
rect 23900 7284 23906 7336
rect 24136 7333 24164 7500
rect 26237 7497 26249 7500
rect 26283 7497 26295 7531
rect 26237 7491 26295 7497
rect 24228 7364 24992 7392
rect 24228 7333 24256 7364
rect 24121 7327 24179 7333
rect 24121 7293 24133 7327
rect 24167 7293 24179 7327
rect 24121 7287 24179 7293
rect 24213 7327 24271 7333
rect 24213 7293 24225 7327
rect 24259 7293 24271 7327
rect 24854 7324 24860 7336
rect 24815 7296 24860 7324
rect 24213 7287 24271 7293
rect 24026 7256 24032 7268
rect 23987 7228 24032 7256
rect 24026 7216 24032 7228
rect 24084 7216 24090 7268
rect 24228 7188 24256 7287
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 24964 7324 24992 7364
rect 25590 7324 25596 7336
rect 24964 7296 25596 7324
rect 25590 7284 25596 7296
rect 25648 7284 25654 7336
rect 25102 7259 25160 7265
rect 25102 7256 25114 7259
rect 24412 7228 25114 7256
rect 24412 7197 24440 7228
rect 25102 7225 25114 7228
rect 25148 7225 25160 7259
rect 25102 7219 25160 7225
rect 23676 7160 24256 7188
rect 24397 7191 24455 7197
rect 24397 7157 24409 7191
rect 24443 7157 24455 7191
rect 24397 7151 24455 7157
rect 1104 7098 28428 7120
rect 1104 7046 10090 7098
rect 10142 7046 10154 7098
rect 10206 7046 10218 7098
rect 10270 7046 10282 7098
rect 10334 7046 19198 7098
rect 19250 7046 19262 7098
rect 19314 7046 19326 7098
rect 19378 7046 19390 7098
rect 19442 7046 28428 7098
rect 1104 7024 28428 7046
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4120 6956 4568 6984
rect 4120 6944 4126 6956
rect 2032 6919 2090 6925
rect 2032 6885 2044 6919
rect 2078 6916 2090 6919
rect 2682 6916 2688 6928
rect 2078 6888 2688 6916
rect 2078 6885 2090 6888
rect 2032 6879 2090 6885
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 4540 6925 4568 6956
rect 7208 6956 7788 6984
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6885 4583 6919
rect 5721 6919 5779 6925
rect 5721 6916 5733 6919
rect 4525 6879 4583 6885
rect 4724 6888 5733 6916
rect 4724 6860 4752 6888
rect 5721 6885 5733 6888
rect 5767 6885 5779 6919
rect 5721 6879 5779 6885
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 2464 6820 2820 6848
rect 2464 6808 2470 6820
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 1780 6644 1808 6743
rect 2792 6712 2820 6820
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4433 6851 4491 6857
rect 4304 6820 4349 6848
rect 4304 6808 4310 6820
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 4706 6848 4712 6860
rect 4663 6820 4712 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4448 6780 4476 6811
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 6178 6848 6184 6860
rect 5583 6820 6040 6848
rect 6139 6820 6184 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 5350 6780 5356 6792
rect 4448 6752 5356 6780
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 4246 6712 4252 6724
rect 2792 6684 4252 6712
rect 4246 6672 4252 6684
rect 4304 6672 4310 6724
rect 6012 6712 6040 6820
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 7208 6848 7236 6956
rect 7650 6916 7656 6928
rect 7484 6888 7656 6916
rect 7374 6848 7380 6860
rect 6696 6820 7236 6848
rect 7335 6820 7380 6848
rect 6696 6808 6702 6820
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 7484 6857 7512 6888
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 7760 6916 7788 6956
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 11388 6956 11437 6984
rect 11388 6944 11394 6956
rect 11425 6953 11437 6956
rect 11471 6953 11483 6987
rect 11425 6947 11483 6953
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 23842 6984 23848 6996
rect 18564 6956 23848 6984
rect 18564 6944 18570 6956
rect 23842 6944 23848 6956
rect 23900 6944 23906 6996
rect 24854 6944 24860 6996
rect 24912 6984 24918 6996
rect 26050 6984 26056 6996
rect 24912 6956 26056 6984
rect 24912 6944 24918 6956
rect 26050 6944 26056 6956
rect 26108 6944 26114 6996
rect 11146 6916 11152 6928
rect 7760 6888 7880 6916
rect 11107 6888 11152 6916
rect 7469 6851 7527 6857
rect 7469 6817 7481 6851
rect 7515 6817 7527 6851
rect 7742 6848 7748 6860
rect 7703 6820 7748 6848
rect 7469 6811 7527 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 7852 6848 7880 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 17586 6916 17592 6928
rect 15764 6888 17592 6916
rect 10870 6848 10876 6860
rect 7852 6820 10456 6848
rect 10831 6820 10876 6848
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 9674 6780 9680 6792
rect 7239 6752 9680 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 7282 6712 7288 6724
rect 6012 6684 7288 6712
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 7653 6715 7711 6721
rect 7653 6681 7665 6715
rect 7699 6712 7711 6715
rect 8110 6712 8116 6724
rect 7699 6684 8116 6712
rect 7699 6681 7711 6684
rect 7653 6675 7711 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 10428 6712 10456 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11054 6848 11060 6860
rect 11015 6820 11060 6848
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12434 6848 12440 6860
rect 12207 6820 12440 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10686 6780 10692 6792
rect 10560 6752 10692 6780
rect 10560 6740 10566 6752
rect 10686 6740 10692 6752
rect 10744 6780 10750 6792
rect 11256 6780 11284 6811
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 15764 6857 15792 6888
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 20254 6916 20260 6928
rect 17880 6888 18184 6916
rect 20215 6888 20260 6916
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6817 15807 6851
rect 15749 6811 15807 6817
rect 16016 6851 16074 6857
rect 16016 6817 16028 6851
rect 16062 6848 16074 6851
rect 16390 6848 16396 6860
rect 16062 6820 16396 6848
rect 16062 6817 16074 6820
rect 16016 6811 16074 6817
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17880 6848 17908 6888
rect 18046 6848 18052 6860
rect 17000 6820 17908 6848
rect 18007 6820 18052 6848
rect 17000 6808 17006 6820
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18156 6848 18184 6888
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 21008 6888 21312 6916
rect 18693 6851 18751 6857
rect 18693 6848 18705 6851
rect 18156 6820 18705 6848
rect 18693 6817 18705 6820
rect 18739 6817 18751 6851
rect 18693 6811 18751 6817
rect 18782 6808 18788 6860
rect 18840 6808 18846 6860
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 20809 6851 20867 6857
rect 20809 6817 20821 6851
rect 20855 6848 20867 6851
rect 21008 6848 21036 6888
rect 21082 6857 21088 6860
rect 20855 6820 21036 6848
rect 20855 6817 20867 6820
rect 20809 6811 20867 6817
rect 21076 6811 21088 6857
rect 21140 6848 21146 6860
rect 21284 6848 21312 6888
rect 22462 6876 22468 6928
rect 22520 6916 22526 6928
rect 22894 6919 22952 6925
rect 22894 6916 22906 6919
rect 22520 6888 22906 6916
rect 22520 6876 22526 6888
rect 22894 6885 22906 6888
rect 22940 6885 22952 6919
rect 23860 6916 23888 6944
rect 25130 6916 25136 6928
rect 23860 6888 25136 6916
rect 22894 6879 22952 6885
rect 25130 6876 25136 6888
rect 25188 6916 25194 6928
rect 25498 6916 25504 6928
rect 25188 6888 25268 6916
rect 25459 6888 25504 6916
rect 25188 6876 25194 6888
rect 21140 6820 21176 6848
rect 21284 6820 22094 6848
rect 11790 6780 11796 6792
rect 10744 6752 11796 6780
rect 10744 6740 10750 6752
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 18800 6780 18828 6808
rect 18187 6752 18828 6780
rect 20180 6780 20208 6811
rect 21082 6808 21088 6811
rect 21140 6808 21146 6820
rect 22066 6780 22094 6820
rect 23198 6808 23204 6860
rect 23256 6848 23262 6860
rect 24578 6848 24584 6860
rect 23256 6820 24584 6848
rect 23256 6808 23262 6820
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 25240 6857 25268 6888
rect 25498 6876 25504 6888
rect 25556 6916 25562 6928
rect 25556 6888 26648 6916
rect 25556 6876 25562 6888
rect 25225 6851 25283 6857
rect 25225 6817 25237 6851
rect 25271 6817 25283 6851
rect 25406 6848 25412 6860
rect 25367 6820 25412 6848
rect 25225 6811 25283 6817
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 25590 6848 25596 6860
rect 25551 6820 25596 6848
rect 25590 6808 25596 6820
rect 25648 6808 25654 6860
rect 26493 6851 26551 6857
rect 26493 6848 26505 6851
rect 25792 6820 26505 6848
rect 22462 6780 22468 6792
rect 20180 6752 20852 6780
rect 22066 6752 22468 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 11882 6712 11888 6724
rect 10428 6684 11888 6712
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 17862 6672 17868 6724
rect 17920 6712 17926 6724
rect 18785 6715 18843 6721
rect 18785 6712 18797 6715
rect 17920 6684 18797 6712
rect 17920 6672 17926 6684
rect 18785 6681 18797 6684
rect 18831 6681 18843 6715
rect 18785 6675 18843 6681
rect 20824 6656 20852 6752
rect 22462 6740 22468 6752
rect 22520 6780 22526 6792
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 22520 6752 22661 6780
rect 22520 6740 22526 6752
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 23658 6672 23664 6724
rect 23716 6712 23722 6724
rect 25792 6721 25820 6820
rect 26493 6817 26505 6820
rect 26539 6817 26551 6851
rect 26620 6848 26648 6888
rect 26620 6820 27660 6848
rect 26493 6811 26551 6817
rect 26050 6740 26056 6792
rect 26108 6780 26114 6792
rect 26237 6783 26295 6789
rect 26237 6780 26249 6783
rect 26108 6752 26249 6780
rect 26108 6740 26114 6752
rect 26237 6749 26249 6752
rect 26283 6749 26295 6783
rect 26237 6743 26295 6749
rect 27632 6721 27660 6820
rect 25777 6715 25835 6721
rect 23716 6684 24164 6712
rect 23716 6672 23722 6684
rect 2130 6644 2136 6656
rect 1780 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 3142 6644 3148 6656
rect 3103 6616 3148 6644
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 3476 6616 4813 6644
rect 3476 6604 3482 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 4801 6607 4859 6613
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7466 6644 7472 6656
rect 7064 6616 7472 6644
rect 7064 6604 7070 6616
rect 7466 6604 7472 6616
rect 7524 6644 7530 6656
rect 10134 6644 10140 6656
rect 7524 6616 10140 6644
rect 7524 6604 7530 6616
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6644 12311 6647
rect 12986 6644 12992 6656
rect 12299 6616 12992 6644
rect 12299 6613 12311 6616
rect 12253 6607 12311 6613
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16540 6616 17141 6644
rect 16540 6604 16546 6616
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 22189 6647 22247 6653
rect 22189 6644 22201 6647
rect 20864 6616 22201 6644
rect 20864 6604 20870 6616
rect 22189 6613 22201 6616
rect 22235 6613 22247 6647
rect 22189 6607 22247 6613
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 24029 6647 24087 6653
rect 24029 6644 24041 6647
rect 22888 6616 24041 6644
rect 22888 6604 22894 6616
rect 24029 6613 24041 6616
rect 24075 6613 24087 6647
rect 24136 6644 24164 6684
rect 25777 6681 25789 6715
rect 25823 6681 25835 6715
rect 25777 6675 25835 6681
rect 27617 6715 27675 6721
rect 27617 6681 27629 6715
rect 27663 6681 27675 6715
rect 27617 6675 27675 6681
rect 26878 6644 26884 6656
rect 24136 6616 26884 6644
rect 24029 6607 24087 6613
rect 26878 6604 26884 6616
rect 26936 6604 26942 6656
rect 1104 6554 28428 6576
rect 1104 6502 5536 6554
rect 5588 6502 5600 6554
rect 5652 6502 5664 6554
rect 5716 6502 5728 6554
rect 5780 6502 14644 6554
rect 14696 6502 14708 6554
rect 14760 6502 14772 6554
rect 14824 6502 14836 6554
rect 14888 6502 23752 6554
rect 23804 6502 23816 6554
rect 23868 6502 23880 6554
rect 23932 6502 23944 6554
rect 23996 6502 28428 6554
rect 1104 6480 28428 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 3234 6440 3240 6452
rect 1627 6412 3240 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 4120 6412 4261 6440
rect 4120 6400 4126 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 6638 6440 6644 6452
rect 5675 6412 6644 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8168 6412 8401 6440
rect 8168 6400 8174 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 8389 6403 8447 6409
rect 9401 6443 9459 6449
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 10778 6440 10784 6452
rect 9447 6412 10784 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 10778 6400 10784 6412
rect 10836 6440 10842 6452
rect 13081 6443 13139 6449
rect 13081 6440 13093 6443
rect 10836 6412 13093 6440
rect 10836 6400 10842 6412
rect 13081 6409 13093 6412
rect 13127 6409 13139 6443
rect 16390 6440 16396 6452
rect 16351 6412 16396 6440
rect 13081 6403 13139 6409
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17678 6440 17684 6452
rect 17639 6412 17684 6440
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 21082 6440 21088 6452
rect 21043 6412 21088 6440
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 23566 6440 23572 6452
rect 22066 6412 23572 6440
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 22066 6372 22094 6412
rect 23566 6400 23572 6412
rect 23624 6400 23630 6452
rect 23845 6443 23903 6449
rect 23845 6409 23857 6443
rect 23891 6440 23903 6443
rect 24302 6440 24308 6452
rect 23891 6412 24308 6440
rect 23891 6409 23903 6412
rect 23845 6403 23903 6409
rect 24302 6400 24308 6412
rect 24360 6400 24366 6452
rect 24397 6443 24455 6449
rect 24397 6409 24409 6443
rect 24443 6409 24455 6443
rect 24397 6403 24455 6409
rect 5408 6344 22094 6372
rect 5408 6332 5414 6344
rect 22830 6332 22836 6384
rect 22888 6372 22894 6384
rect 24412 6372 24440 6403
rect 24578 6400 24584 6452
rect 24636 6440 24642 6452
rect 26789 6443 26847 6449
rect 26789 6440 26801 6443
rect 24636 6412 26801 6440
rect 24636 6400 24642 6412
rect 26789 6409 26801 6412
rect 26835 6409 26847 6443
rect 26789 6403 26847 6409
rect 22888 6344 24440 6372
rect 22888 6332 22894 6344
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4304 6276 4997 6304
rect 4304 6264 4310 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12308 6276 12725 6304
rect 12308 6264 12314 6276
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 19337 6307 19395 6313
rect 17368 6276 18920 6304
rect 17368 6264 17374 6276
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 3136 6239 3194 6245
rect 3136 6205 3148 6239
rect 3182 6236 3194 6239
rect 3418 6236 3424 6248
rect 3182 6208 3424 6236
rect 3182 6205 3194 6208
rect 3136 6199 3194 6205
rect 2130 6128 2136 6180
rect 2188 6168 2194 6180
rect 2884 6168 2912 6199
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 4847 6208 5457 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5445 6205 5457 6208
rect 5491 6236 5503 6239
rect 7006 6236 7012 6248
rect 5491 6208 7012 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8096 6239 8154 6245
rect 8096 6236 8108 6239
rect 7708 6208 8108 6236
rect 7708 6196 7714 6208
rect 8096 6205 8108 6208
rect 8142 6205 8154 6239
rect 8096 6199 8154 6205
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 8478 6236 8484 6248
rect 8439 6208 8484 6236
rect 8205 6199 8263 6205
rect 4062 6168 4068 6180
rect 2188 6140 4068 6168
rect 2188 6128 2194 6140
rect 4062 6128 4068 6140
rect 4120 6128 4126 6180
rect 8220 6168 8248 6199
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8588 6208 8953 6236
rect 8386 6168 8392 6180
rect 8220 6140 8392 6168
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8588 6100 8616 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 9122 6236 9128 6248
rect 9083 6208 9128 6236
rect 8941 6199 8999 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9493 6239 9551 6245
rect 9272 6208 9317 6236
rect 9272 6196 9278 6208
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 10502 6236 10508 6248
rect 9539 6208 10508 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 12618 6236 12624 6248
rect 12579 6208 12624 6236
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12802 6236 12808 6248
rect 12763 6208 12808 6236
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13173 6239 13231 6245
rect 12952 6208 12997 6236
rect 12952 6196 12958 6208
rect 13173 6205 13185 6239
rect 13219 6205 13231 6239
rect 13998 6236 14004 6248
rect 13959 6208 14004 6236
rect 13173 6199 13231 6205
rect 7975 6072 8616 6100
rect 8941 6103 8999 6109
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9490 6100 9496 6112
rect 8987 6072 9496 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 13188 6100 13216 6199
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14182 6236 14188 6248
rect 14143 6208 14188 6236
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 14366 6236 14372 6248
rect 14327 6208 14372 6236
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 15194 6196 15200 6248
rect 15252 6236 15258 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 15252 6208 15393 6236
rect 15252 6196 15258 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 15838 6236 15844 6248
rect 15799 6208 15844 6236
rect 15381 6199 15439 6205
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6236 16267 6239
rect 16390 6236 16396 6248
rect 16255 6208 16396 6236
rect 16255 6205 16267 6208
rect 16209 6199 16267 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 17402 6196 17408 6248
rect 17460 6236 17466 6248
rect 17497 6239 17555 6245
rect 17497 6236 17509 6239
rect 17460 6208 17509 6236
rect 17460 6196 17466 6208
rect 17497 6205 17509 6208
rect 17543 6236 17555 6239
rect 17862 6236 17868 6248
rect 17543 6208 17868 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 17862 6196 17868 6208
rect 17920 6236 17926 6248
rect 18325 6239 18383 6245
rect 18325 6236 18337 6239
rect 17920 6208 18337 6236
rect 17920 6196 17926 6208
rect 18325 6205 18337 6208
rect 18371 6205 18383 6239
rect 18892 6236 18920 6276
rect 19337 6273 19349 6307
rect 19383 6304 19395 6307
rect 19383 6276 20944 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 20530 6236 20536 6248
rect 18892 6208 19288 6236
rect 20491 6208 20536 6236
rect 18325 6199 18383 6205
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14277 6171 14335 6177
rect 14277 6168 14289 6171
rect 13780 6140 14289 6168
rect 13780 6128 13786 6140
rect 14277 6137 14289 6140
rect 14323 6137 14335 6171
rect 14277 6131 14335 6137
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 16025 6171 16083 6177
rect 16025 6168 16037 6171
rect 14700 6140 16037 6168
rect 14700 6128 14706 6140
rect 16025 6137 16037 6140
rect 16071 6137 16083 6171
rect 16025 6131 16083 6137
rect 16117 6171 16175 6177
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 16482 6168 16488 6180
rect 16163 6140 16488 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 16482 6128 16488 6140
rect 16540 6128 16546 6180
rect 16942 6128 16948 6180
rect 17000 6168 17006 6180
rect 19153 6171 19211 6177
rect 19153 6168 19165 6171
rect 17000 6140 19165 6168
rect 17000 6128 17006 6140
rect 19153 6137 19165 6140
rect 19199 6137 19211 6171
rect 19260 6168 19288 6208
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 20806 6236 20812 6248
rect 20767 6208 20812 6236
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 20916 6245 20944 6276
rect 22922 6264 22928 6316
rect 22980 6304 22986 6316
rect 23385 6307 23443 6313
rect 23385 6304 23397 6307
rect 22980 6276 23397 6304
rect 22980 6264 22986 6276
rect 23385 6273 23397 6276
rect 23431 6273 23443 6307
rect 23385 6267 23443 6273
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6236 20959 6239
rect 21266 6236 21272 6248
rect 20947 6208 21272 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 23106 6236 23112 6248
rect 23067 6208 23112 6236
rect 23106 6196 23112 6208
rect 23164 6196 23170 6248
rect 23293 6239 23351 6245
rect 23293 6205 23305 6239
rect 23339 6205 23351 6239
rect 23293 6199 23351 6205
rect 23477 6239 23535 6245
rect 23477 6205 23489 6239
rect 23523 6236 23535 6239
rect 23566 6236 23572 6248
rect 23523 6208 23572 6236
rect 23523 6205 23535 6208
rect 23477 6199 23535 6205
rect 20717 6171 20775 6177
rect 20717 6168 20729 6171
rect 19260 6140 20729 6168
rect 19153 6131 19211 6137
rect 20717 6137 20729 6140
rect 20763 6137 20775 6171
rect 20717 6131 20775 6137
rect 23308 6112 23336 6199
rect 23566 6196 23572 6208
rect 23624 6196 23630 6248
rect 23661 6239 23719 6245
rect 23661 6205 23673 6239
rect 23707 6205 23719 6239
rect 24302 6236 24308 6248
rect 24263 6208 24308 6236
rect 23661 6199 23719 6205
rect 23676 6168 23704 6199
rect 24302 6196 24308 6208
rect 24360 6196 24366 6248
rect 26142 6196 26148 6248
rect 26200 6236 26206 6248
rect 26697 6239 26755 6245
rect 26697 6236 26709 6239
rect 26200 6208 26709 6236
rect 26200 6196 26206 6208
rect 26697 6205 26709 6208
rect 26743 6205 26755 6239
rect 26697 6199 26755 6205
rect 25314 6168 25320 6180
rect 23676 6140 25320 6168
rect 25314 6128 25320 6140
rect 25372 6128 25378 6180
rect 14458 6100 14464 6112
rect 13188 6072 14464 6100
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 15010 6100 15016 6112
rect 14599 6072 15016 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15930 6100 15936 6112
rect 15243 6072 15936 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 16908 6072 18429 6100
rect 16908 6060 16914 6072
rect 18417 6069 18429 6072
rect 18463 6100 18475 6103
rect 22094 6100 22100 6112
rect 18463 6072 22100 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 22094 6060 22100 6072
rect 22152 6060 22158 6112
rect 23290 6060 23296 6112
rect 23348 6060 23354 6112
rect 23658 6060 23664 6112
rect 23716 6100 23722 6112
rect 24670 6100 24676 6112
rect 23716 6072 24676 6100
rect 23716 6060 23722 6072
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 24762 6060 24768 6112
rect 24820 6100 24826 6112
rect 24820 6072 24865 6100
rect 24820 6060 24826 6072
rect 1104 6010 28428 6032
rect 1104 5958 10090 6010
rect 10142 5958 10154 6010
rect 10206 5958 10218 6010
rect 10270 5958 10282 6010
rect 10334 5958 19198 6010
rect 19250 5958 19262 6010
rect 19314 5958 19326 6010
rect 19378 5958 19390 6010
rect 19442 5958 28428 6010
rect 1104 5936 28428 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 5902 5896 5908 5908
rect 4387 5868 5908 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8570 5896 8576 5908
rect 7892 5868 8576 5896
rect 7892 5856 7898 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9916 5868 10057 5896
rect 9916 5856 9922 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 10045 5859 10103 5865
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 10597 5899 10655 5905
rect 10597 5896 10609 5899
rect 10560 5868 10609 5896
rect 10560 5856 10566 5868
rect 10597 5865 10609 5868
rect 10643 5865 10655 5899
rect 10597 5859 10655 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12676 5868 12817 5896
rect 12676 5856 12682 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 12952 5868 14841 5896
rect 12952 5856 12958 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 16574 5856 16580 5908
rect 16632 5896 16638 5908
rect 16853 5899 16911 5905
rect 16853 5896 16865 5899
rect 16632 5868 16865 5896
rect 16632 5856 16638 5868
rect 16853 5865 16865 5868
rect 16899 5865 16911 5899
rect 21545 5899 21603 5905
rect 16853 5859 16911 5865
rect 16960 5868 20668 5896
rect 7460 5831 7518 5837
rect 7460 5797 7472 5831
rect 7506 5828 7518 5831
rect 9769 5831 9827 5837
rect 7506 5800 8524 5828
rect 7506 5797 7518 5800
rect 7460 5791 7518 5797
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 3200 5732 4261 5760
rect 3200 5720 3206 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 8294 5760 8300 5772
rect 7239 5732 8300 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8496 5692 8524 5800
rect 9769 5797 9781 5831
rect 9815 5828 9827 5831
rect 10410 5828 10416 5840
rect 9815 5800 10416 5828
rect 9815 5797 9827 5800
rect 9769 5791 9827 5797
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 13814 5828 13820 5840
rect 13096 5800 13820 5828
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9582 5692 9588 5704
rect 8496 5664 9588 5692
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9692 5692 9720 5723
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 10502 5760 10508 5772
rect 9916 5732 9961 5760
rect 10463 5732 10508 5760
rect 9916 5720 9922 5732
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 10870 5720 10876 5772
rect 10928 5760 10934 5772
rect 11241 5763 11299 5769
rect 11241 5760 11253 5763
rect 10928 5732 11253 5760
rect 10928 5720 10934 5732
rect 11241 5729 11253 5732
rect 11287 5729 11299 5763
rect 11422 5760 11428 5772
rect 11383 5732 11428 5760
rect 11241 5723 11299 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11655 5763 11713 5769
rect 11655 5729 11667 5763
rect 11701 5760 11713 5763
rect 11790 5760 11796 5772
rect 11701 5732 11796 5760
rect 11701 5729 11713 5732
rect 11655 5723 11713 5729
rect 9950 5692 9956 5704
rect 9692 5664 9956 5692
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 11532 5692 11560 5723
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 12986 5760 12992 5772
rect 12947 5732 12992 5760
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13096 5769 13124 5800
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 15102 5828 15108 5840
rect 14752 5800 15108 5828
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13998 5760 14004 5772
rect 13403 5732 14004 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13998 5720 14004 5732
rect 14056 5720 14062 5772
rect 14752 5769 14780 5800
rect 15102 5788 15108 5800
rect 15160 5828 15166 5840
rect 16960 5828 16988 5868
rect 15160 5800 16988 5828
rect 15160 5788 15166 5800
rect 17402 5788 17408 5840
rect 17460 5828 17466 5840
rect 18877 5831 18935 5837
rect 18877 5828 18889 5831
rect 17460 5800 18889 5828
rect 17460 5788 17466 5800
rect 18877 5797 18889 5800
rect 18923 5797 18935 5831
rect 18877 5791 18935 5797
rect 19061 5831 19119 5837
rect 19061 5797 19073 5831
rect 19107 5828 19119 5831
rect 20530 5828 20536 5840
rect 19107 5800 20536 5828
rect 19107 5797 19119 5800
rect 19061 5791 19119 5797
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 20640 5828 20668 5868
rect 21545 5865 21557 5899
rect 21591 5896 21603 5899
rect 22554 5896 22560 5908
rect 21591 5868 22560 5896
rect 21591 5865 21603 5868
rect 21545 5859 21603 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 22738 5856 22744 5908
rect 22796 5896 22802 5908
rect 23017 5899 23075 5905
rect 23017 5896 23029 5899
rect 22796 5868 23029 5896
rect 22796 5856 22802 5868
rect 23017 5865 23029 5868
rect 23063 5865 23075 5899
rect 23017 5859 23075 5865
rect 23382 5856 23388 5908
rect 23440 5896 23446 5908
rect 24854 5896 24860 5908
rect 23440 5868 24860 5896
rect 23440 5856 23446 5868
rect 24854 5856 24860 5868
rect 24912 5856 24918 5908
rect 23753 5831 23811 5837
rect 23753 5828 23765 5831
rect 20640 5800 22094 5828
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 15740 5763 15798 5769
rect 15740 5729 15752 5763
rect 15786 5760 15798 5763
rect 16206 5760 16212 5772
rect 15786 5732 16212 5760
rect 15786 5729 15798 5732
rect 15740 5723 15798 5729
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 17000 5732 17509 5760
rect 17000 5720 17006 5732
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 19794 5720 19800 5772
rect 19852 5760 19858 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19852 5732 20177 5760
rect 19852 5720 19858 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 20496 5732 21097 5760
rect 20496 5720 20502 5732
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 21085 5723 21143 5729
rect 12434 5692 12440 5704
rect 11532 5664 12440 5692
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 15473 5695 15531 5701
rect 15473 5692 15485 5695
rect 15344 5664 15485 5692
rect 15344 5652 15350 5664
rect 15473 5661 15485 5664
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 16540 5664 17785 5692
rect 16540 5652 16546 5664
rect 17773 5661 17785 5664
rect 17819 5692 17831 5695
rect 18414 5692 18420 5704
rect 17819 5664 18420 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 14642 5624 14648 5636
rect 2746 5596 4476 5624
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2746 5556 2774 5596
rect 1912 5528 2774 5556
rect 4448 5556 4476 5596
rect 8128 5596 14648 5624
rect 8128 5556 8156 5596
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 22066 5624 22094 5800
rect 22572 5800 23765 5828
rect 22572 5769 22600 5800
rect 23753 5797 23765 5800
rect 23799 5828 23811 5831
rect 24394 5828 24400 5840
rect 23799 5800 24400 5828
rect 23799 5797 23811 5800
rect 23753 5791 23811 5797
rect 24394 5788 24400 5800
rect 24452 5788 24458 5840
rect 27430 5788 27436 5840
rect 27488 5828 27494 5840
rect 27525 5831 27583 5837
rect 27525 5828 27537 5831
rect 27488 5800 27537 5828
rect 27488 5788 27494 5800
rect 27525 5797 27537 5800
rect 27571 5797 27583 5831
rect 27706 5828 27712 5840
rect 27667 5800 27712 5828
rect 27525 5791 27583 5797
rect 27706 5788 27712 5800
rect 27764 5788 27770 5840
rect 22557 5763 22615 5769
rect 22557 5729 22569 5763
rect 22603 5729 22615 5763
rect 22557 5723 22615 5729
rect 22738 5720 22744 5772
rect 22796 5760 22802 5772
rect 23477 5763 23535 5769
rect 23477 5760 23489 5763
rect 22796 5732 23489 5760
rect 22796 5720 22802 5732
rect 23477 5729 23489 5732
rect 23523 5729 23535 5763
rect 23658 5760 23664 5772
rect 23619 5732 23664 5760
rect 23477 5723 23535 5729
rect 23658 5720 23664 5732
rect 23716 5720 23722 5772
rect 23845 5763 23903 5769
rect 23845 5729 23857 5763
rect 23891 5729 23903 5763
rect 23845 5723 23903 5729
rect 23014 5652 23020 5704
rect 23072 5692 23078 5704
rect 23860 5692 23888 5723
rect 23072 5664 23888 5692
rect 23072 5652 23078 5664
rect 27154 5624 27160 5636
rect 19536 5596 21220 5624
rect 22066 5596 27160 5624
rect 4448 5528 8156 5556
rect 1912 5516 1918 5528
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10870 5556 10876 5568
rect 9732 5528 10876 5556
rect 9732 5516 9738 5528
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 11790 5556 11796 5568
rect 11751 5528 11796 5556
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 19536 5556 19564 5596
rect 17276 5528 19564 5556
rect 17276 5516 17282 5528
rect 19610 5516 19616 5568
rect 19668 5556 19674 5568
rect 21192 5565 21220 5596
rect 27154 5584 27160 5596
rect 27212 5584 27218 5636
rect 19981 5559 20039 5565
rect 19981 5556 19993 5559
rect 19668 5528 19993 5556
rect 19668 5516 19674 5528
rect 19981 5525 19993 5528
rect 20027 5525 20039 5559
rect 19981 5519 20039 5525
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 22830 5556 22836 5568
rect 21223 5528 22836 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 24029 5559 24087 5565
rect 24029 5525 24041 5559
rect 24075 5556 24087 5559
rect 24118 5556 24124 5568
rect 24075 5528 24124 5556
rect 24075 5525 24087 5528
rect 24029 5519 24087 5525
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 1104 5466 28428 5488
rect 1104 5414 5536 5466
rect 5588 5414 5600 5466
rect 5652 5414 5664 5466
rect 5716 5414 5728 5466
rect 5780 5414 14644 5466
rect 14696 5414 14708 5466
rect 14760 5414 14772 5466
rect 14824 5414 14836 5466
rect 14888 5414 23752 5466
rect 23804 5414 23816 5466
rect 23868 5414 23880 5466
rect 23932 5414 23944 5466
rect 23996 5414 28428 5466
rect 1104 5392 28428 5414
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 3878 5352 3884 5364
rect 3559 5324 3884 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 7742 5352 7748 5364
rect 7239 5324 7748 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 7742 5312 7748 5324
rect 7800 5312 7806 5364
rect 22278 5352 22284 5364
rect 10888 5324 22284 5352
rect 7650 5244 7656 5296
rect 7708 5284 7714 5296
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7708 5256 7849 5284
rect 7708 5244 7714 5256
rect 7837 5253 7849 5256
rect 7883 5253 7895 5287
rect 7837 5247 7895 5253
rect 9490 5244 9496 5296
rect 9548 5284 9554 5296
rect 10781 5287 10839 5293
rect 10781 5284 10793 5287
rect 9548 5256 10793 5284
rect 9548 5244 9554 5256
rect 10781 5253 10793 5256
rect 10827 5253 10839 5287
rect 10781 5247 10839 5253
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8352 5188 8401 5216
rect 8352 5176 8358 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 10888 5216 10916 5324
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 22830 5352 22836 5364
rect 22520 5324 22836 5352
rect 22520 5312 22526 5324
rect 22830 5312 22836 5324
rect 22888 5352 22894 5364
rect 23382 5352 23388 5364
rect 22888 5324 23388 5352
rect 22888 5312 22894 5324
rect 23382 5312 23388 5324
rect 23440 5352 23446 5364
rect 23440 5324 23796 5352
rect 23440 5312 23446 5324
rect 12526 5284 12532 5296
rect 9824 5188 10916 5216
rect 11532 5256 12532 5284
rect 9824 5176 9830 5188
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 10428 5157 10456 5188
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 10229 5151 10287 5157
rect 10229 5117 10241 5151
rect 10275 5117 10287 5151
rect 10229 5111 10287 5117
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5148 10655 5151
rect 11532 5148 11560 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 14458 5244 14464 5296
rect 14516 5284 14522 5296
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 14516 5256 15117 5284
rect 14516 5244 14522 5256
rect 15105 5253 15117 5256
rect 15151 5253 15163 5287
rect 15105 5247 15163 5253
rect 16206 5244 16212 5296
rect 16264 5284 16270 5296
rect 16393 5287 16451 5293
rect 16393 5284 16405 5287
rect 16264 5256 16405 5284
rect 16264 5244 16270 5256
rect 16393 5253 16405 5256
rect 16439 5253 16451 5287
rect 16393 5247 16451 5253
rect 17678 5244 17684 5296
rect 17736 5284 17742 5296
rect 21542 5284 21548 5296
rect 17736 5256 19104 5284
rect 21503 5256 21548 5284
rect 17736 5244 17742 5256
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 14148 5188 15148 5216
rect 14148 5176 14154 5188
rect 12066 5148 12072 5160
rect 10643 5120 11560 5148
rect 12027 5120 12072 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 2400 5083 2458 5089
rect 2400 5049 2412 5083
rect 2446 5080 2458 5083
rect 2774 5080 2780 5092
rect 2446 5052 2780 5080
rect 2446 5049 2458 5052
rect 2400 5043 2458 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 7760 5012 7788 5111
rect 8656 5083 8714 5089
rect 8656 5049 8668 5083
rect 8702 5080 8714 5083
rect 9950 5080 9956 5092
rect 8702 5052 9956 5080
rect 8702 5049 8714 5052
rect 8656 5043 8714 5049
rect 9950 5040 9956 5052
rect 10008 5040 10014 5092
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 7760 4984 9781 5012
rect 9769 4981 9781 4984
rect 9815 5012 9827 5015
rect 9858 5012 9864 5024
rect 9815 4984 9864 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10244 5012 10272 5111
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12526 5148 12532 5160
rect 12483 5120 12532 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 13078 5148 13084 5160
rect 12860 5120 13084 5148
rect 12860 5108 12866 5120
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14292 5120 15025 5148
rect 10502 5040 10508 5092
rect 10560 5080 10566 5092
rect 10560 5052 10605 5080
rect 10560 5040 10566 5052
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 12250 5080 12256 5092
rect 11480 5052 12256 5080
rect 11480 5040 11486 5052
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 12345 5083 12403 5089
rect 12345 5049 12357 5083
rect 12391 5080 12403 5083
rect 13348 5083 13406 5089
rect 12391 5052 13308 5080
rect 12391 5049 12403 5052
rect 12345 5043 12403 5049
rect 12066 5012 12072 5024
rect 10244 4984 12072 5012
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 13280 5012 13308 5052
rect 13348 5049 13360 5083
rect 13394 5080 13406 5083
rect 13446 5080 13452 5092
rect 13394 5052 13452 5080
rect 13394 5049 13406 5052
rect 13348 5043 13406 5049
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 13538 5012 13544 5024
rect 13280 4984 13544 5012
rect 13538 4972 13544 4984
rect 13596 5012 13602 5024
rect 14292 5012 14320 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 15120 5080 15148 5188
rect 15856 5188 17601 5216
rect 15856 5160 15884 5188
rect 17589 5185 17601 5188
rect 17635 5216 17647 5219
rect 17954 5216 17960 5228
rect 17635 5188 17960 5216
rect 17635 5185 17647 5188
rect 17589 5179 17647 5185
rect 17954 5176 17960 5188
rect 18012 5216 18018 5228
rect 18012 5188 18092 5216
rect 18012 5176 18018 5188
rect 15838 5148 15844 5160
rect 15799 5120 15844 5148
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16209 5151 16267 5157
rect 16209 5117 16221 5151
rect 16255 5148 16267 5151
rect 16482 5148 16488 5160
rect 16255 5120 16488 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 17402 5148 17408 5160
rect 17363 5120 17408 5148
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 18064 5157 18092 5188
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 19076 5225 19104 5256
rect 21542 5244 21548 5256
rect 21600 5244 21606 5296
rect 23768 5225 23796 5324
rect 24394 5312 24400 5364
rect 24452 5352 24458 5364
rect 25133 5355 25191 5361
rect 25133 5352 25145 5355
rect 24452 5324 25145 5352
rect 24452 5312 24458 5324
rect 25133 5321 25145 5324
rect 25179 5321 25191 5355
rect 25133 5315 25191 5321
rect 19061 5219 19119 5225
rect 18196 5188 18828 5216
rect 18196 5176 18202 5188
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18414 5148 18420 5160
rect 18327 5120 18420 5148
rect 18049 5111 18107 5117
rect 18414 5108 18420 5120
rect 18472 5148 18478 5160
rect 18690 5148 18696 5160
rect 18472 5120 18696 5148
rect 18472 5108 18478 5120
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 18800 5148 18828 5188
rect 19061 5185 19073 5219
rect 19107 5185 19119 5219
rect 23753 5219 23811 5225
rect 19061 5179 19119 5185
rect 22066 5188 22968 5216
rect 20990 5148 20996 5160
rect 18800 5120 20996 5148
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21453 5151 21511 5157
rect 21453 5117 21465 5151
rect 21499 5148 21511 5151
rect 22066 5148 22094 5188
rect 22940 5160 22968 5188
rect 23753 5185 23765 5219
rect 23799 5185 23811 5219
rect 27614 5216 27620 5228
rect 23753 5179 23811 5185
rect 24780 5188 27620 5216
rect 22649 5151 22707 5157
rect 22649 5148 22661 5151
rect 21499 5120 22094 5148
rect 22204 5120 22661 5148
rect 21499 5117 21511 5120
rect 21453 5111 21511 5117
rect 16025 5083 16083 5089
rect 16025 5080 16037 5083
rect 15120 5052 16037 5080
rect 16025 5049 16037 5052
rect 16071 5049 16083 5083
rect 16025 5043 16083 5049
rect 16117 5083 16175 5089
rect 16117 5049 16129 5083
rect 16163 5080 16175 5083
rect 16574 5080 16580 5092
rect 16163 5052 16580 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 18230 5080 18236 5092
rect 18191 5052 18236 5080
rect 18230 5040 18236 5052
rect 18288 5040 18294 5092
rect 18325 5083 18383 5089
rect 18325 5049 18337 5083
rect 18371 5080 18383 5083
rect 19328 5083 19386 5089
rect 18371 5052 19288 5080
rect 18371 5049 18383 5052
rect 18325 5043 18383 5049
rect 14458 5012 14464 5024
rect 13596 4984 14320 5012
rect 14371 4984 14464 5012
rect 13596 4972 13602 4984
rect 14458 4972 14464 4984
rect 14516 5012 14522 5024
rect 15102 5012 15108 5024
rect 14516 4984 15108 5012
rect 14516 4972 14522 4984
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 18601 5015 18659 5021
rect 18601 4981 18613 5015
rect 18647 5012 18659 5015
rect 19058 5012 19064 5024
rect 18647 4984 19064 5012
rect 18647 4981 18659 4984
rect 18601 4975 18659 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 19260 5012 19288 5052
rect 19328 5049 19340 5083
rect 19374 5080 19386 5083
rect 19518 5080 19524 5092
rect 19374 5052 19524 5080
rect 19374 5049 19386 5052
rect 19328 5043 19386 5049
rect 19518 5040 19524 5052
rect 19576 5040 19582 5092
rect 22094 5040 22100 5092
rect 22152 5080 22158 5092
rect 22204 5080 22232 5120
rect 22649 5117 22661 5120
rect 22695 5148 22707 5151
rect 22738 5148 22744 5160
rect 22695 5120 22744 5148
rect 22695 5117 22707 5120
rect 22649 5111 22707 5117
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 22922 5148 22928 5160
rect 22883 5120 22928 5148
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 23014 5108 23020 5160
rect 23072 5148 23078 5160
rect 24780 5148 24808 5188
rect 27614 5176 27620 5188
rect 27672 5176 27678 5228
rect 23072 5120 23117 5148
rect 23676 5120 24808 5148
rect 26697 5151 26755 5157
rect 23072 5108 23078 5120
rect 22152 5052 22232 5080
rect 22152 5040 22158 5052
rect 22370 5040 22376 5092
rect 22428 5080 22434 5092
rect 22833 5083 22891 5089
rect 22833 5080 22845 5083
rect 22428 5052 22845 5080
rect 22428 5040 22434 5052
rect 22833 5049 22845 5052
rect 22879 5049 22891 5083
rect 23676 5080 23704 5120
rect 26697 5117 26709 5151
rect 26743 5148 26755 5151
rect 26878 5148 26884 5160
rect 26743 5120 26884 5148
rect 26743 5117 26755 5120
rect 26697 5111 26755 5117
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 22833 5043 22891 5049
rect 23032 5052 23704 5080
rect 24020 5083 24078 5089
rect 19978 5012 19984 5024
rect 19260 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20438 5012 20444 5024
rect 20399 4984 20444 5012
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 23032 5012 23060 5052
rect 24020 5049 24032 5083
rect 24066 5080 24078 5083
rect 24118 5080 24124 5092
rect 24066 5052 24124 5080
rect 24066 5049 24078 5052
rect 24020 5043 24078 5049
rect 24118 5040 24124 5052
rect 24176 5040 24182 5092
rect 23198 5012 23204 5024
rect 22336 4984 23060 5012
rect 23159 4984 23204 5012
rect 22336 4972 22342 4984
rect 23198 4972 23204 4984
rect 23256 4972 23262 5024
rect 24394 4972 24400 5024
rect 24452 5012 24458 5024
rect 26881 5015 26939 5021
rect 26881 5012 26893 5015
rect 24452 4984 26893 5012
rect 24452 4972 24458 4984
rect 26881 4981 26893 4984
rect 26927 4981 26939 5015
rect 26881 4975 26939 4981
rect 1104 4922 28428 4944
rect 1104 4870 10090 4922
rect 10142 4870 10154 4922
rect 10206 4870 10218 4922
rect 10270 4870 10282 4922
rect 10334 4870 19198 4922
rect 19250 4870 19262 4922
rect 19314 4870 19326 4922
rect 19378 4870 19390 4922
rect 19442 4870 28428 4922
rect 1104 4848 28428 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 6825 4811 6883 4817
rect 1636 4780 6132 4808
rect 1636 4768 1642 4780
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 1762 4740 1768 4752
rect 1719 4712 1768 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 1762 4700 1768 4712
rect 1820 4700 1826 4752
rect 2406 4740 2412 4752
rect 2332 4712 2412 4740
rect 2332 4681 2360 4712
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 3878 4740 3884 4752
rect 2639 4712 3884 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4641 2375 4675
rect 2498 4672 2504 4684
rect 2459 4644 2504 4672
rect 2317 4635 2375 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 2866 4672 2872 4684
rect 2731 4644 2872 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 4890 4632 4896 4684
rect 4948 4672 4954 4684
rect 5057 4675 5115 4681
rect 5057 4672 5069 4675
rect 4948 4644 5069 4672
rect 4948 4632 4954 4644
rect 5057 4641 5069 4644
rect 5103 4641 5115 4675
rect 5057 4635 5115 4641
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4798 4604 4804 4616
rect 4212 4576 4804 4604
rect 4212 4564 4218 4576
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 6104 4604 6132 4780
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 6914 4808 6920 4820
rect 6871 4780 6920 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 9122 4808 9128 4820
rect 8527 4780 9128 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 10008 4780 10149 4808
rect 10008 4768 10014 4780
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10137 4771 10195 4777
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 13446 4808 13452 4820
rect 13407 4780 13452 4808
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 20533 4811 20591 4817
rect 14844 4780 20484 4808
rect 9674 4740 9680 4752
rect 9600 4712 9680 4740
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6236 4644 6745 4672
rect 6236 4632 6242 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 8478 4672 8484 4684
rect 8435 4644 8484 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 9600 4681 9628 4712
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9824 4712 9869 4740
rect 9824 4700 9830 4712
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9858 4672 9864 4684
rect 9819 4644 9864 4672
rect 9585 4635 9643 4641
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10704 4672 10732 4768
rect 11324 4743 11382 4749
rect 11324 4709 11336 4743
rect 11370 4740 11382 4743
rect 11790 4740 11796 4752
rect 11370 4712 11796 4740
rect 11370 4709 11382 4712
rect 11324 4703 11382 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 12250 4700 12256 4752
rect 12308 4740 12314 4752
rect 13081 4743 13139 4749
rect 13081 4740 13093 4743
rect 12308 4712 13093 4740
rect 12308 4700 12314 4712
rect 13081 4709 13093 4712
rect 13127 4740 13139 4743
rect 14844 4740 14872 4780
rect 15010 4749 15016 4752
rect 15004 4740 15016 4749
rect 13127 4712 14872 4740
rect 14971 4712 15016 4740
rect 13127 4709 13139 4712
rect 13081 4703 13139 4709
rect 15004 4703 15016 4712
rect 15010 4700 15016 4703
rect 15068 4700 15074 4752
rect 16942 4700 16948 4752
rect 17000 4740 17006 4752
rect 17037 4743 17095 4749
rect 17037 4740 17049 4743
rect 17000 4712 17049 4740
rect 17000 4700 17006 4712
rect 17037 4709 17049 4712
rect 17083 4709 17095 4743
rect 17037 4703 17095 4709
rect 17948 4743 18006 4749
rect 17948 4709 17960 4743
rect 17994 4740 18006 4743
rect 19702 4740 19708 4752
rect 17994 4712 19708 4740
rect 17994 4709 18006 4712
rect 17948 4703 18006 4709
rect 19702 4700 19708 4712
rect 19760 4700 19766 4752
rect 20254 4700 20260 4752
rect 20312 4740 20318 4752
rect 20456 4740 20484 4780
rect 20533 4777 20545 4811
rect 20579 4808 20591 4811
rect 20622 4808 20628 4820
rect 20579 4780 20628 4808
rect 20579 4777 20591 4780
rect 20533 4771 20591 4777
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 20990 4808 20996 4820
rect 20951 4780 20996 4808
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 22922 4768 22928 4820
rect 22980 4808 22986 4820
rect 24213 4811 24271 4817
rect 24213 4808 24225 4811
rect 22980 4780 24225 4808
rect 22980 4768 22986 4780
rect 24213 4777 24225 4780
rect 24259 4777 24271 4811
rect 24213 4771 24271 4777
rect 23100 4743 23158 4749
rect 20312 4712 20357 4740
rect 20456 4712 21947 4740
rect 20312 4700 20318 4712
rect 9999 4644 10732 4672
rect 11057 4675 11115 4681
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 12802 4672 12808 4684
rect 11103 4644 12808 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4641 12955 4675
rect 12897 4635 12955 4641
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4641 13231 4675
rect 13173 4635 13231 4641
rect 6104 4576 9674 4604
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 2869 4539 2927 4545
rect 2869 4536 2881 4539
rect 2832 4508 2881 4536
rect 2832 4496 2838 4508
rect 2869 4505 2881 4508
rect 2915 4505 2927 4539
rect 2869 4499 2927 4505
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4468 1823 4471
rect 2958 4468 2964 4480
rect 1811 4440 2964 4468
rect 1811 4437 1823 4440
rect 1765 4431 1823 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 6178 4468 6184 4480
rect 6139 4440 6184 4468
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 9646 4468 9674 4576
rect 12158 4564 12164 4616
rect 12216 4604 12222 4616
rect 12912 4604 12940 4635
rect 12216 4576 12940 4604
rect 12216 4564 12222 4576
rect 13188 4536 13216 4635
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 14737 4675 14795 4681
rect 13320 4644 13365 4672
rect 13320 4632 13326 4644
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15286 4672 15292 4684
rect 14783 4644 15292 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 17678 4672 17684 4684
rect 17639 4644 17684 4672
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 17770 4632 17776 4684
rect 17828 4672 17834 4684
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 17828 4644 19993 4672
rect 17828 4632 17834 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 20162 4672 20168 4684
rect 20123 4644 20168 4672
rect 19981 4635 20039 4641
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 20349 4675 20407 4681
rect 20349 4641 20361 4675
rect 20395 4641 20407 4675
rect 21174 4672 21180 4684
rect 21135 4644 21180 4672
rect 20349 4635 20407 4641
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 20364 4604 20392 4635
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4641 21879 4675
rect 21919 4672 21947 4712
rect 23100 4709 23112 4743
rect 23146 4740 23158 4743
rect 23198 4740 23204 4752
rect 23146 4712 23204 4740
rect 23146 4709 23158 4712
rect 23100 4703 23158 4709
rect 23198 4700 23204 4712
rect 23256 4700 23262 4752
rect 27522 4740 27528 4752
rect 27483 4712 27528 4740
rect 27522 4700 27528 4712
rect 27580 4700 27586 4752
rect 25406 4672 25412 4684
rect 21919 4644 23888 4672
rect 25367 4644 25412 4672
rect 21821 4635 21879 4641
rect 18748 4576 20392 4604
rect 18748 4564 18754 4576
rect 14458 4536 14464 4548
rect 13188 4508 14464 4536
rect 14458 4496 14464 4508
rect 14516 4496 14522 4548
rect 17218 4536 17224 4548
rect 17179 4508 17224 4536
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 18966 4496 18972 4548
rect 19024 4536 19030 4548
rect 21637 4539 21695 4545
rect 21637 4536 21649 4539
rect 19024 4508 21649 4536
rect 19024 4496 19030 4508
rect 21637 4505 21649 4508
rect 21683 4505 21695 4539
rect 21637 4499 21695 4505
rect 14090 4468 14096 4480
rect 9646 4440 14096 4468
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 14366 4428 14372 4480
rect 14424 4468 14430 4480
rect 16117 4471 16175 4477
rect 16117 4468 16129 4471
rect 14424 4440 16129 4468
rect 14424 4428 14430 4440
rect 16117 4437 16129 4440
rect 16163 4437 16175 4471
rect 16117 4431 16175 4437
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 18104 4440 19073 4468
rect 18104 4428 18110 4440
rect 19061 4437 19073 4440
rect 19107 4468 19119 4471
rect 20254 4468 20260 4480
rect 19107 4440 20260 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 20346 4428 20352 4480
rect 20404 4468 20410 4480
rect 21836 4468 21864 4635
rect 22830 4604 22836 4616
rect 22791 4576 22836 4604
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 23860 4604 23888 4644
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 26050 4632 26056 4684
rect 26108 4672 26114 4684
rect 26145 4675 26203 4681
rect 26145 4672 26157 4675
rect 26108 4644 26157 4672
rect 26108 4632 26114 4644
rect 26145 4641 26157 4644
rect 26191 4641 26203 4675
rect 26786 4672 26792 4684
rect 26747 4644 26792 4672
rect 26145 4635 26203 4641
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 27709 4607 27767 4613
rect 27709 4604 27721 4607
rect 23860 4576 27721 4604
rect 27709 4573 27721 4576
rect 27755 4573 27767 4607
rect 27709 4567 27767 4573
rect 24210 4496 24216 4548
rect 24268 4536 24274 4548
rect 26973 4539 27031 4545
rect 26973 4536 26985 4539
rect 24268 4508 26985 4536
rect 24268 4496 24274 4508
rect 26973 4505 26985 4508
rect 27019 4505 27031 4539
rect 26973 4499 27031 4505
rect 25222 4468 25228 4480
rect 20404 4440 21864 4468
rect 25183 4440 25228 4468
rect 20404 4428 20410 4440
rect 25222 4428 25228 4440
rect 25280 4428 25286 4480
rect 26326 4468 26332 4480
rect 26287 4440 26332 4468
rect 26326 4428 26332 4440
rect 26384 4428 26390 4480
rect 1104 4378 28428 4400
rect 1104 4326 5536 4378
rect 5588 4326 5600 4378
rect 5652 4326 5664 4378
rect 5716 4326 5728 4378
rect 5780 4326 14644 4378
rect 14696 4326 14708 4378
rect 14760 4326 14772 4378
rect 14824 4326 14836 4378
rect 14888 4326 23752 4378
rect 23804 4326 23816 4378
rect 23868 4326 23880 4378
rect 23932 4326 23944 4378
rect 23996 4326 28428 4378
rect 1104 4304 28428 4326
rect 2498 4264 2504 4276
rect 2459 4236 2504 4264
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 10321 4267 10379 4273
rect 10321 4233 10333 4267
rect 10367 4264 10379 4267
rect 10502 4264 10508 4276
rect 10367 4236 10508 4264
rect 10367 4233 10379 4236
rect 10321 4227 10379 4233
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 12434 4264 12440 4276
rect 12084 4236 12440 4264
rect 6178 4128 6184 4140
rect 4632 4100 6184 4128
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 2774 4060 2780 4072
rect 2731 4032 2780 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 3142 4060 3148 4072
rect 3103 4032 3148 4060
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 4632 4069 4660 4100
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8352 4100 8953 4128
rect 8352 4088 8358 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 12084 4137 12112 4236
rect 12434 4224 12440 4236
rect 12492 4264 12498 4276
rect 12802 4264 12808 4276
rect 12492 4236 12808 4264
rect 12492 4224 12498 4236
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 13538 4264 13544 4276
rect 13495 4236 13544 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 14645 4267 14703 4273
rect 14645 4264 14657 4267
rect 13648 4236 14657 4264
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 13648 4196 13676 4236
rect 14645 4233 14657 4236
rect 14691 4233 14703 4267
rect 14645 4227 14703 4233
rect 18230 4224 18236 4276
rect 18288 4264 18294 4276
rect 26326 4264 26332 4276
rect 18288 4236 26332 4264
rect 18288 4224 18294 4236
rect 26326 4224 26332 4236
rect 26384 4224 26390 4276
rect 13412 4168 13676 4196
rect 13832 4168 14136 4196
rect 13412 4156 13418 4168
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10468 4100 11069 4128
rect 10468 4088 10474 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13832 4128 13860 4168
rect 13998 4128 14004 4140
rect 13136 4100 13860 4128
rect 13959 4100 14004 4128
rect 13136 4088 13142 4100
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14108 4128 14136 4168
rect 15286 4156 15292 4208
rect 15344 4196 15350 4208
rect 17678 4196 17684 4208
rect 15344 4168 17684 4196
rect 15344 4156 15350 4168
rect 17678 4156 17684 4168
rect 17736 4196 17742 4208
rect 17736 4168 18276 4196
rect 17736 4156 17742 4168
rect 18138 4128 18144 4140
rect 14108 4100 18144 4128
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18248 4128 18276 4168
rect 18322 4156 18328 4208
rect 18380 4196 18386 4208
rect 18966 4196 18972 4208
rect 18380 4168 18972 4196
rect 18380 4156 18386 4168
rect 18966 4156 18972 4168
rect 19024 4156 19030 4208
rect 19978 4156 19984 4208
rect 20036 4196 20042 4208
rect 20349 4199 20407 4205
rect 20349 4196 20361 4199
rect 20036 4168 20361 4196
rect 20036 4156 20042 4168
rect 20349 4165 20361 4168
rect 20395 4165 20407 4199
rect 20349 4159 20407 4165
rect 18414 4128 18420 4140
rect 18248 4100 18420 4128
rect 18414 4088 18420 4100
rect 18472 4128 18478 4140
rect 18472 4100 19012 4128
rect 18472 4088 18478 4100
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 4304 4032 4353 4060
rect 4304 4020 4310 4032
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 2866 3992 2872 4004
rect 1903 3964 2872 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1452 3896 1961 3924
rect 1452 3884 1458 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 3329 3927 3387 3933
rect 3329 3924 3341 3927
rect 2648 3896 3341 3924
rect 2648 3884 2654 3896
rect 3329 3893 3341 3896
rect 3375 3893 3387 3927
rect 4356 3924 4384 4023
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 5350 4060 5356 4072
rect 4764 4032 4809 4060
rect 5311 4032 5356 4060
rect 4764 4020 4770 4032
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5460 4032 5733 4060
rect 4522 3992 4528 4004
rect 4483 3964 4528 3992
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 4724 3992 4752 4020
rect 5460 3992 5488 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 9208 4063 9266 4069
rect 9208 4029 9220 4063
rect 9254 4060 9266 4063
rect 9490 4060 9496 4072
rect 9254 4032 9496 4060
rect 9254 4029 9266 4032
rect 9208 4023 9266 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 12158 4060 12164 4072
rect 9876 4032 12164 4060
rect 9876 4004 9904 4032
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 12336 4063 12394 4069
rect 12336 4029 12348 4063
rect 12382 4060 12394 4063
rect 12618 4060 12624 4072
rect 12382 4032 12624 4060
rect 12382 4029 12394 4032
rect 12336 4023 12394 4029
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 13906 4060 13912 4072
rect 13867 4032 13912 4060
rect 13906 4020 13912 4032
rect 13964 4020 13970 4072
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14148 4032 14565 4060
rect 14148 4020 14154 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 14553 4023 14611 4029
rect 14640 4032 15209 4060
rect 4724 3964 5488 3992
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3961 5595 3995
rect 5537 3955 5595 3961
rect 5629 3995 5687 4001
rect 5629 3961 5641 3995
rect 5675 3992 5687 3995
rect 7098 3992 7104 4004
rect 5675 3964 7104 3992
rect 5675 3961 5687 3964
rect 5629 3955 5687 3961
rect 5350 3924 5356 3936
rect 4356 3896 5356 3924
rect 3329 3887 3387 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5552 3924 5580 3955
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 9674 3992 9680 4004
rect 7248 3964 9680 3992
rect 7248 3952 7254 3964
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 9858 3952 9864 4004
rect 9916 3952 9922 4004
rect 10873 3995 10931 4001
rect 10873 3961 10885 3995
rect 10919 3992 10931 3995
rect 12526 3992 12532 4004
rect 10919 3964 12532 3992
rect 10919 3961 10931 3964
rect 10873 3955 10931 3961
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 14640 3992 14668 4032
rect 15197 4029 15209 4032
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 17000 4032 17325 4060
rect 17000 4020 17006 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17954 4060 17960 4072
rect 17915 4032 17960 4060
rect 17313 4023 17371 4029
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4060 18383 4063
rect 18690 4060 18696 4072
rect 18371 4032 18696 4060
rect 18371 4029 18383 4032
rect 18325 4023 18383 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 18984 4069 19012 4100
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21634 4128 21640 4140
rect 20772 4100 21640 4128
rect 20772 4088 20778 4100
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 22646 4128 22652 4140
rect 22607 4100 22652 4128
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 23290 4128 23296 4140
rect 23251 4100 23296 4128
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 18969 4063 19027 4069
rect 18969 4029 18981 4063
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 19058 4020 19064 4072
rect 19116 4060 19122 4072
rect 19225 4063 19283 4069
rect 19225 4060 19237 4063
rect 19116 4032 19237 4060
rect 19116 4020 19122 4032
rect 19225 4029 19237 4032
rect 19271 4029 19283 4063
rect 19225 4023 19283 4029
rect 21082 4020 21088 4072
rect 21140 4060 21146 4072
rect 21177 4063 21235 4069
rect 21177 4060 21189 4063
rect 21140 4032 21189 4060
rect 21140 4020 21146 4032
rect 21177 4029 21189 4032
rect 21223 4029 21235 4063
rect 21177 4023 21235 4029
rect 22002 4020 22008 4072
rect 22060 4060 22066 4072
rect 22557 4063 22615 4069
rect 22557 4060 22569 4063
rect 22060 4032 22569 4060
rect 22060 4020 22066 4032
rect 22557 4029 22569 4032
rect 22603 4029 22615 4063
rect 23198 4060 23204 4072
rect 23159 4032 23204 4060
rect 22557 4023 22615 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23382 4020 23388 4072
rect 23440 4060 23446 4072
rect 24029 4063 24087 4069
rect 24029 4060 24041 4063
rect 23440 4032 24041 4060
rect 23440 4020 23446 4032
rect 24029 4029 24041 4032
rect 24075 4029 24087 4063
rect 24854 4060 24860 4072
rect 24815 4032 24860 4060
rect 24029 4023 24087 4029
rect 24854 4020 24860 4032
rect 24912 4020 24918 4072
rect 25958 4060 25964 4072
rect 25919 4032 25964 4060
rect 25958 4020 25964 4032
rect 26016 4020 26022 4072
rect 13412 3964 14668 3992
rect 13412 3952 13418 3964
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 16209 3995 16267 4001
rect 16209 3992 16221 3995
rect 15160 3964 16221 3992
rect 15160 3952 15166 3964
rect 16209 3961 16221 3964
rect 16255 3961 16267 3995
rect 16209 3955 16267 3961
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 17405 3995 17463 4001
rect 17405 3992 17417 3995
rect 16724 3964 17417 3992
rect 16724 3952 16730 3964
rect 17405 3961 17417 3964
rect 17451 3961 17463 3995
rect 17405 3955 17463 3961
rect 18141 3995 18199 4001
rect 18141 3961 18153 3995
rect 18187 3961 18199 3995
rect 18141 3955 18199 3961
rect 5718 3924 5724 3936
rect 5552 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 12986 3924 12992 3936
rect 7984 3896 12992 3924
rect 7984 3884 7990 3896
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 14090 3924 14096 3936
rect 13228 3896 14096 3924
rect 13228 3884 13234 3896
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 16172 3896 16313 3924
rect 16172 3884 16178 3896
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 18156 3924 18184 3955
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18288 3964 18333 3992
rect 22112 3964 23888 3992
rect 18288 3952 18294 3964
rect 18322 3924 18328 3936
rect 18156 3896 18328 3924
rect 16301 3887 16359 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3924 18567 3927
rect 19518 3924 19524 3936
rect 18555 3896 19524 3924
rect 18555 3893 18567 3896
rect 18509 3887 18567 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 22112 3924 22140 3964
rect 20220 3896 22140 3924
rect 20220 3884 20226 3896
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 23382 3924 23388 3936
rect 22704 3896 23388 3924
rect 22704 3884 22710 3896
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 23860 3933 23888 3964
rect 23934 3952 23940 4004
rect 23992 3992 23998 4004
rect 26697 3995 26755 4001
rect 26697 3992 26709 3995
rect 23992 3964 26709 3992
rect 23992 3952 23998 3964
rect 26697 3961 26709 3964
rect 26743 3961 26755 3995
rect 26697 3955 26755 3961
rect 26881 3995 26939 4001
rect 26881 3961 26893 3995
rect 26927 3992 26939 3995
rect 27614 3992 27620 4004
rect 26927 3964 27620 3992
rect 26927 3961 26939 3964
rect 26881 3955 26939 3961
rect 27614 3952 27620 3964
rect 27672 3952 27678 4004
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 24946 3884 24952 3936
rect 25004 3924 25010 3936
rect 25041 3927 25099 3933
rect 25041 3924 25053 3927
rect 25004 3896 25053 3924
rect 25004 3884 25010 3896
rect 25041 3893 25053 3896
rect 25087 3893 25099 3927
rect 26142 3924 26148 3936
rect 26103 3896 26148 3924
rect 25041 3887 25099 3893
rect 26142 3884 26148 3896
rect 26200 3884 26206 3936
rect 1104 3834 28428 3856
rect 1104 3782 10090 3834
rect 10142 3782 10154 3834
rect 10206 3782 10218 3834
rect 10270 3782 10282 3834
rect 10334 3782 19198 3834
rect 19250 3782 19262 3834
rect 19314 3782 19326 3834
rect 19378 3782 19390 3834
rect 19442 3782 28428 3834
rect 1104 3760 28428 3782
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 6917 3723 6975 3729
rect 5776 3692 6868 3720
rect 5776 3680 5782 3692
rect 5804 3655 5862 3661
rect 5804 3621 5816 3655
rect 5850 3652 5862 3655
rect 5902 3652 5908 3664
rect 5850 3624 5908 3652
rect 5850 3621 5862 3624
rect 5804 3615 5862 3621
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 6840 3652 6868 3692
rect 6917 3689 6929 3723
rect 6963 3720 6975 3723
rect 7098 3720 7104 3732
rect 6963 3692 7104 3720
rect 6963 3689 6975 3692
rect 6917 3683 6975 3689
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 8956 3692 12848 3720
rect 8956 3652 8984 3692
rect 6840 3624 8984 3652
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 10229 3655 10287 3661
rect 10229 3652 10241 3655
rect 9640 3624 10241 3652
rect 9640 3612 9646 3624
rect 10229 3621 10241 3624
rect 10275 3621 10287 3655
rect 12434 3652 12440 3664
rect 10229 3615 10287 3621
rect 10980 3624 12440 3652
rect 1486 3584 1492 3596
rect 1447 3556 1492 3584
rect 1486 3544 1492 3556
rect 1544 3544 1550 3596
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 1820 3556 2145 3584
rect 1820 3544 1826 3556
rect 2133 3553 2145 3556
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2372 3556 2881 3584
rect 2372 3544 2378 3556
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 5537 3587 5595 3593
rect 5537 3584 5549 3587
rect 4856 3556 5549 3584
rect 4856 3544 4862 3556
rect 5537 3553 5549 3556
rect 5583 3553 5595 3587
rect 5537 3547 5595 3553
rect 7834 3544 7840 3596
rect 7892 3584 7898 3596
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 7892 3556 7941 3584
rect 7892 3544 7898 3556
rect 7929 3553 7941 3556
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8754 3584 8760 3596
rect 8435 3556 8760 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9916 3556 9965 3584
rect 9916 3544 9922 3556
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10686 3584 10692 3596
rect 10367 3556 10692 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 9674 3516 9680 3528
rect 8720 3488 9680 3516
rect 8720 3476 8726 3488
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 10152 3516 10180 3547
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10980 3593 11008 3624
rect 12434 3612 12440 3624
rect 12492 3612 12498 3664
rect 12820 3652 12848 3692
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 18969 3723 19027 3729
rect 18969 3720 18981 3723
rect 12952 3692 18981 3720
rect 12952 3680 12958 3692
rect 18969 3689 18981 3692
rect 19015 3689 19027 3723
rect 18969 3683 19027 3689
rect 19702 3680 19708 3732
rect 19760 3720 19766 3732
rect 21174 3720 21180 3732
rect 19760 3692 21180 3720
rect 19760 3680 19766 3692
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 23014 3680 23020 3732
rect 23072 3720 23078 3732
rect 23842 3720 23848 3732
rect 23072 3692 23848 3720
rect 23072 3680 23078 3692
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 13081 3655 13139 3661
rect 12820 3624 12940 3652
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 11232 3587 11290 3593
rect 11232 3553 11244 3587
rect 11278 3584 11290 3587
rect 12710 3584 12716 3596
rect 11278 3556 12716 3584
rect 11278 3553 11290 3556
rect 11232 3547 11290 3553
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 9824 3488 10180 3516
rect 9824 3476 9830 3488
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12820 3516 12848 3547
rect 12032 3488 12848 3516
rect 12912 3516 12940 3624
rect 13081 3621 13093 3655
rect 13127 3652 13139 3655
rect 13906 3652 13912 3664
rect 13127 3624 13912 3652
rect 13127 3621 13139 3624
rect 13081 3615 13139 3621
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 14366 3612 14372 3664
rect 14424 3652 14430 3664
rect 14921 3655 14979 3661
rect 14921 3652 14933 3655
rect 14424 3624 14933 3652
rect 14424 3612 14430 3624
rect 14921 3621 14933 3624
rect 14967 3621 14979 3655
rect 14921 3615 14979 3621
rect 15028 3624 16896 3652
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 13173 3587 13231 3593
rect 13044 3556 13089 3584
rect 13044 3544 13050 3556
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 13262 3584 13268 3596
rect 13219 3556 13268 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 15028 3516 15056 3624
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15654 3584 15660 3596
rect 15151 3556 15660 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 15832 3587 15890 3593
rect 15832 3553 15844 3587
rect 15878 3584 15890 3587
rect 16758 3584 16764 3596
rect 15878 3556 16764 3584
rect 15878 3553 15890 3556
rect 15832 3547 15890 3553
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 12912 3488 15056 3516
rect 12032 3476 12038 3488
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15344 3488 15577 3516
rect 15344 3476 15350 3488
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 16868 3516 16896 3624
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 20438 3652 20444 3664
rect 18288 3624 20444 3652
rect 18288 3612 18294 3624
rect 20438 3612 20444 3624
rect 20496 3612 20502 3664
rect 20901 3655 20959 3661
rect 20901 3621 20913 3655
rect 20947 3652 20959 3655
rect 22002 3652 22008 3664
rect 20947 3624 22008 3652
rect 20947 3621 20959 3624
rect 20901 3615 20959 3621
rect 22002 3612 22008 3624
rect 22060 3612 22066 3664
rect 22738 3612 22744 3664
rect 22796 3652 22802 3664
rect 23661 3655 23719 3661
rect 22796 3624 23520 3652
rect 22796 3612 22802 3624
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17405 3587 17463 3593
rect 17405 3584 17417 3587
rect 17092 3556 17417 3584
rect 17092 3544 17098 3556
rect 17405 3553 17417 3556
rect 17451 3553 17463 3587
rect 17405 3547 17463 3553
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 18141 3587 18199 3593
rect 18141 3584 18153 3587
rect 18104 3556 18153 3584
rect 18104 3544 18110 3556
rect 18141 3553 18153 3556
rect 18187 3553 18199 3587
rect 18874 3584 18880 3596
rect 18835 3556 18880 3584
rect 18141 3547 18199 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 19978 3584 19984 3596
rect 19939 3556 19984 3584
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20530 3544 20536 3596
rect 20588 3584 20594 3596
rect 20625 3587 20683 3593
rect 20625 3584 20637 3587
rect 20588 3556 20637 3584
rect 20588 3544 20594 3556
rect 20625 3553 20637 3556
rect 20671 3553 20683 3587
rect 20625 3547 20683 3553
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 20993 3587 21051 3593
rect 20993 3553 21005 3587
rect 21039 3584 21051 3587
rect 21266 3584 21272 3596
rect 21039 3556 21272 3584
rect 21039 3553 21051 3556
rect 20993 3547 21051 3553
rect 20254 3516 20260 3528
rect 16868 3488 20260 3516
rect 15565 3479 15623 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20824 3516 20852 3547
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 21904 3587 21962 3593
rect 21904 3553 21916 3587
rect 21950 3584 21962 3587
rect 23382 3584 23388 3596
rect 21950 3556 23388 3584
rect 21950 3553 21962 3556
rect 21904 3547 21962 3553
rect 23382 3544 23388 3556
rect 23440 3544 23446 3596
rect 23492 3593 23520 3624
rect 23661 3621 23673 3655
rect 23707 3652 23719 3655
rect 25222 3652 25228 3664
rect 23707 3624 25228 3652
rect 23707 3621 23719 3624
rect 23661 3615 23719 3621
rect 25222 3612 25228 3624
rect 25280 3612 25286 3664
rect 25593 3655 25651 3661
rect 25593 3621 25605 3655
rect 25639 3652 25651 3655
rect 25682 3652 25688 3664
rect 25639 3624 25688 3652
rect 25639 3621 25651 3624
rect 25593 3615 25651 3621
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 26329 3655 26387 3661
rect 26329 3621 26341 3655
rect 26375 3652 26387 3655
rect 26510 3652 26516 3664
rect 26375 3624 26516 3652
rect 26375 3621 26387 3624
rect 26329 3615 26387 3621
rect 26510 3612 26516 3624
rect 26568 3612 26574 3664
rect 23477 3587 23535 3593
rect 23477 3553 23489 3587
rect 23523 3553 23535 3587
rect 23477 3547 23535 3553
rect 23753 3587 23811 3593
rect 23753 3553 23765 3587
rect 23799 3553 23811 3587
rect 23753 3547 23811 3553
rect 20364 3488 20852 3516
rect 21637 3519 21695 3525
rect 7745 3451 7803 3457
rect 7745 3417 7757 3451
rect 7791 3448 7803 3451
rect 9490 3448 9496 3460
rect 7791 3420 9496 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 12345 3451 12403 3457
rect 9600 3420 10640 3448
rect 934 3340 940 3392
rect 992 3380 998 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 992 3352 1593 3380
rect 992 3340 998 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 4062 3380 4068 3392
rect 3099 3352 4068 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 6604 3352 8585 3380
rect 6604 3340 6610 3352
rect 8573 3349 8585 3352
rect 8619 3349 8631 3383
rect 8573 3343 8631 3349
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9600 3380 9628 3420
rect 10502 3380 10508 3392
rect 8720 3352 9628 3380
rect 10463 3352 10508 3380
rect 8720 3340 8726 3352
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 10612 3380 10640 3420
rect 12345 3417 12357 3451
rect 12391 3448 12403 3451
rect 12526 3448 12532 3460
rect 12391 3420 12532 3448
rect 12391 3417 12403 3420
rect 12345 3411 12403 3417
rect 12526 3408 12532 3420
rect 12584 3448 12590 3460
rect 13170 3448 13176 3460
rect 12584 3420 13176 3448
rect 12584 3408 12590 3420
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 15470 3448 15476 3460
rect 13280 3420 15476 3448
rect 13280 3380 13308 3420
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 20364 3448 20392 3488
rect 21637 3485 21649 3519
rect 21683 3485 21695 3519
rect 23768 3516 23796 3547
rect 23842 3544 23848 3596
rect 23900 3584 23906 3596
rect 23900 3556 23945 3584
rect 23900 3544 23906 3556
rect 24394 3544 24400 3596
rect 24452 3584 24458 3596
rect 25406 3584 25412 3596
rect 24452 3556 25412 3584
rect 24452 3544 24458 3556
rect 25406 3544 25412 3556
rect 25464 3544 25470 3596
rect 26418 3544 26424 3596
rect 26476 3584 26482 3596
rect 26973 3587 27031 3593
rect 26973 3584 26985 3587
rect 26476 3556 26985 3584
rect 26476 3544 26482 3556
rect 26973 3553 26985 3556
rect 27019 3584 27031 3587
rect 27062 3584 27068 3596
rect 27019 3556 27068 3584
rect 27019 3553 27031 3556
rect 26973 3547 27031 3553
rect 27062 3544 27068 3556
rect 27120 3544 27126 3596
rect 24302 3516 24308 3528
rect 23768 3488 24308 3516
rect 21637 3479 21695 3485
rect 16500 3420 20392 3448
rect 10612 3352 13308 3380
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 13538 3380 13544 3392
rect 13403 3352 13544 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 16500 3380 16528 3420
rect 20438 3408 20444 3460
rect 20496 3448 20502 3460
rect 21652 3448 21680 3479
rect 24302 3476 24308 3488
rect 24360 3516 24366 3528
rect 24762 3516 24768 3528
rect 24360 3488 24768 3516
rect 24360 3476 24366 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25774 3448 25780 3460
rect 20496 3420 21680 3448
rect 25735 3420 25780 3448
rect 20496 3408 20502 3420
rect 25774 3408 25780 3420
rect 25832 3408 25838 3460
rect 26510 3448 26516 3460
rect 26471 3420 26516 3448
rect 26510 3408 26516 3420
rect 26568 3408 26574 3460
rect 16942 3380 16948 3392
rect 13780 3352 16528 3380
rect 16903 3352 16948 3380
rect 13780 3340 13786 3352
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 18230 3380 18236 3392
rect 18191 3352 18236 3380
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19024 3352 20085 3380
rect 19024 3340 19030 3352
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 21174 3380 21180 3392
rect 21135 3352 21180 3380
rect 20073 3343 20131 3349
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 23017 3383 23075 3389
rect 23017 3349 23029 3383
rect 23063 3380 23075 3383
rect 23198 3380 23204 3392
rect 23063 3352 23204 3380
rect 23063 3349 23075 3352
rect 23017 3343 23075 3349
rect 23198 3340 23204 3352
rect 23256 3340 23262 3392
rect 24029 3383 24087 3389
rect 24029 3349 24041 3383
rect 24075 3380 24087 3383
rect 24118 3380 24124 3392
rect 24075 3352 24124 3380
rect 24075 3349 24087 3352
rect 24029 3343 24087 3349
rect 24118 3340 24124 3352
rect 24176 3340 24182 3392
rect 1104 3290 28428 3312
rect 1104 3238 5536 3290
rect 5588 3238 5600 3290
rect 5652 3238 5664 3290
rect 5716 3238 5728 3290
rect 5780 3238 14644 3290
rect 14696 3238 14708 3290
rect 14760 3238 14772 3290
rect 14824 3238 14836 3290
rect 14888 3238 23752 3290
rect 23804 3238 23816 3290
rect 23868 3238 23880 3290
rect 23932 3238 23944 3290
rect 23996 3238 28428 3290
rect 1104 3216 28428 3238
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4522 3176 4528 3188
rect 4387 3148 4528 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 13722 3176 13728 3188
rect 5215 3148 13728 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 13906 3176 13912 3188
rect 13867 3148 13912 3176
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 18046 3176 18052 3188
rect 16132 3148 18052 3176
rect 1581 3111 1639 3117
rect 1581 3077 1593 3111
rect 1627 3108 1639 3111
rect 1627 3080 8800 3108
rect 1627 3077 1639 3080
rect 1581 3071 1639 3077
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 8662 3040 8668 3052
rect 1544 3012 8668 3040
rect 1544 3000 1550 3012
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 2148 2981 2176 3012
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 8772 3040 8800 3080
rect 9766 3068 9772 3120
rect 9824 3108 9830 3120
rect 12250 3108 12256 3120
rect 9824 3080 12256 3108
rect 9824 3068 9830 3080
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 12434 3068 12440 3120
rect 12492 3108 12498 3120
rect 12492 3080 12572 3108
rect 12492 3068 12498 3080
rect 12342 3040 12348 3052
rect 8772 3012 8892 3040
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2941 2191 2975
rect 2866 2972 2872 2984
rect 2827 2944 2872 2972
rect 2133 2935 2191 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3602 2972 3608 2984
rect 3563 2944 3608 2972
rect 3602 2932 3608 2944
rect 3660 2932 3666 2984
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4525 2975 4583 2981
rect 4525 2972 4537 2975
rect 4212 2944 4537 2972
rect 4212 2932 4218 2944
rect 4525 2941 4537 2944
rect 4571 2941 4583 2975
rect 4525 2935 4583 2941
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2941 5043 2975
rect 6914 2972 6920 2984
rect 6875 2944 6920 2972
rect 4985 2935 5043 2941
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 5000 2904 5028 2935
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 8352 2944 8769 2972
rect 8352 2932 8358 2944
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 3292 2876 5028 2904
rect 8864 2904 8892 3012
rect 10612 3012 12348 3040
rect 9024 2975 9082 2981
rect 9024 2941 9036 2975
rect 9070 2972 9082 2975
rect 10502 2972 10508 2984
rect 9070 2944 10508 2972
rect 9070 2941 9082 2944
rect 9024 2935 9082 2941
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 10612 2904 10640 3012
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12544 3049 12572 3080
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 12434 2972 12440 2984
rect 11011 2944 12440 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 12796 2975 12854 2981
rect 12796 2941 12808 2975
rect 12842 2972 12854 2975
rect 13538 2972 13544 2984
rect 12842 2944 13544 2972
rect 12842 2941 12854 2944
rect 12796 2935 12854 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 13688 2944 14473 2972
rect 13688 2932 13694 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 15102 2972 15108 2984
rect 15015 2944 15108 2972
rect 14461 2935 14519 2941
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15841 2975 15899 2981
rect 15841 2941 15853 2975
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 8864 2876 10640 2904
rect 11149 2907 11207 2913
rect 3292 2864 3298 2876
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 11974 2904 11980 2916
rect 11195 2876 11980 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 12894 2864 12900 2916
rect 12952 2904 12958 2916
rect 15120 2904 15148 2932
rect 12952 2876 15148 2904
rect 15856 2904 15884 2935
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16132 2981 16160 3148
rect 18046 3136 18052 3148
rect 18104 3176 18110 3188
rect 18693 3179 18751 3185
rect 18693 3176 18705 3179
rect 18104 3148 18705 3176
rect 18104 3136 18110 3148
rect 18693 3145 18705 3148
rect 18739 3145 18751 3179
rect 18693 3139 18751 3145
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 21361 3179 21419 3185
rect 21361 3176 21373 3179
rect 19208 3148 21373 3176
rect 19208 3136 19214 3148
rect 21361 3145 21373 3148
rect 21407 3145 21419 3179
rect 21361 3139 21419 3145
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 24820 3148 24869 3176
rect 24820 3136 24826 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 20364 3080 22094 3108
rect 16390 3040 16396 3052
rect 16224 3012 16396 3040
rect 16224 2981 16252 3012
rect 16390 3000 16396 3012
rect 16448 3040 16454 3052
rect 17218 3040 17224 3052
rect 16448 3012 17224 3040
rect 16448 3000 16454 3012
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 18414 3000 18420 3052
rect 18472 3040 18478 3052
rect 19325 3040 19331 3052
rect 19383 3049 19389 3052
rect 18472 3012 19331 3040
rect 18472 3000 18478 3012
rect 19325 3000 19331 3012
rect 19383 3040 19395 3049
rect 19383 3012 19476 3040
rect 19383 3003 19395 3012
rect 19383 3000 19389 3003
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15988 2944 16037 2972
rect 15988 2932 15994 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16025 2935 16083 2941
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 16209 2975 16267 2981
rect 16209 2941 16221 2975
rect 16255 2941 16267 2975
rect 16850 2972 16856 2984
rect 16209 2935 16267 2941
rect 16316 2944 16856 2972
rect 16316 2904 16344 2944
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 18432 2972 18460 3000
rect 19886 2972 19892 2984
rect 17359 2944 18460 2972
rect 19536 2944 19892 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 17558 2907 17616 2913
rect 17558 2904 17570 2907
rect 15856 2876 16344 2904
rect 16408 2876 17570 2904
rect 12952 2864 12958 2876
rect 16040 2848 16068 2876
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 10137 2839 10195 2845
rect 10137 2836 10149 2839
rect 9640 2808 10149 2836
rect 9640 2796 9646 2808
rect 10137 2805 10149 2808
rect 10183 2805 10195 2839
rect 10137 2799 10195 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 12492 2808 14565 2836
rect 12492 2796 12498 2808
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 14553 2799 14611 2805
rect 16022 2796 16028 2848
rect 16080 2796 16086 2848
rect 16408 2845 16436 2876
rect 17558 2873 17570 2876
rect 17604 2873 17616 2907
rect 17558 2867 17616 2873
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 19536 2904 19564 2944
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 20364 2972 20392 3080
rect 20128 2944 20392 2972
rect 20128 2932 20134 2944
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 21269 2975 21327 2981
rect 21269 2972 21281 2975
rect 20772 2944 21281 2972
rect 20772 2932 20778 2944
rect 21269 2941 21281 2944
rect 21315 2941 21327 2975
rect 22066 2972 22094 3080
rect 22830 3000 22836 3052
rect 22888 3040 22894 3052
rect 23477 3043 23535 3049
rect 23477 3040 23489 3043
rect 22888 3012 23489 3040
rect 22888 3000 22894 3012
rect 23477 3009 23489 3012
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 22066 2944 22661 2972
rect 21269 2935 21327 2941
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 23744 2975 23802 2981
rect 23744 2941 23756 2975
rect 23790 2972 23802 2975
rect 24118 2972 24124 2984
rect 23790 2944 24124 2972
rect 23790 2941 23802 2944
rect 23744 2935 23802 2941
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 25314 2932 25320 2984
rect 25372 2972 25378 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25372 2944 25973 2972
rect 25372 2932 25378 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 26697 2975 26755 2981
rect 26697 2941 26709 2975
rect 26743 2972 26755 2975
rect 27338 2972 27344 2984
rect 26743 2944 27344 2972
rect 26743 2941 26755 2944
rect 26697 2935 26755 2941
rect 27338 2932 27344 2944
rect 27396 2932 27402 2984
rect 18288 2876 19564 2904
rect 19604 2907 19662 2913
rect 18288 2864 18294 2876
rect 19604 2873 19616 2907
rect 19650 2904 19662 2907
rect 20162 2904 20168 2916
rect 19650 2876 20168 2904
rect 19650 2873 19662 2876
rect 19604 2867 19662 2873
rect 20162 2864 20168 2876
rect 20220 2864 20226 2916
rect 26145 2907 26203 2913
rect 26145 2873 26157 2907
rect 26191 2904 26203 2907
rect 26234 2904 26240 2916
rect 26191 2876 26240 2904
rect 26191 2873 26203 2876
rect 26145 2867 26203 2873
rect 26234 2864 26240 2876
rect 26292 2864 26298 2916
rect 16393 2839 16451 2845
rect 16393 2805 16405 2839
rect 16439 2805 16451 2839
rect 16393 2799 16451 2805
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 20346 2836 20352 2848
rect 18012 2808 20352 2836
rect 18012 2796 18018 2808
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 20680 2808 20729 2836
rect 20680 2796 20686 2808
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 21634 2796 21640 2848
rect 21692 2836 21698 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 21692 2808 22753 2836
rect 21692 2796 21698 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 22741 2799 22799 2805
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 24762 2836 24768 2848
rect 23532 2808 24768 2836
rect 23532 2796 23538 2808
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 26786 2836 26792 2848
rect 26747 2808 26792 2836
rect 26786 2796 26792 2808
rect 26844 2796 26850 2848
rect 1104 2746 28428 2768
rect 1104 2694 10090 2746
rect 10142 2694 10154 2746
rect 10206 2694 10218 2746
rect 10270 2694 10282 2746
rect 10334 2694 19198 2746
rect 19250 2694 19262 2746
rect 19314 2694 19326 2746
rect 19378 2694 19390 2746
rect 19442 2694 28428 2746
rect 1104 2672 28428 2694
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 5905 2635 5963 2641
rect 3660 2604 5856 2632
rect 3660 2592 3666 2604
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 4798 2564 4804 2576
rect 4571 2536 4804 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 5828 2564 5856 2604
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6454 2632 6460 2644
rect 5951 2604 6460 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 9490 2592 9496 2644
rect 9548 2632 9554 2644
rect 9548 2604 12664 2632
rect 9548 2592 9554 2604
rect 10413 2567 10471 2573
rect 10413 2564 10425 2567
rect 5828 2536 10425 2564
rect 10413 2533 10425 2536
rect 10459 2533 10471 2567
rect 12526 2564 12532 2576
rect 12487 2536 12532 2564
rect 10413 2527 10471 2533
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 12636 2564 12664 2604
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 12768 2604 12817 2632
rect 12768 2592 12774 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 16758 2632 16764 2644
rect 16623 2604 16764 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19383 2604 19748 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 16209 2567 16267 2573
rect 16209 2564 16221 2567
rect 12636 2536 16221 2564
rect 16209 2533 16221 2536
rect 16255 2533 16267 2567
rect 16209 2527 16267 2533
rect 16301 2567 16359 2573
rect 16301 2533 16313 2567
rect 16347 2564 16359 2567
rect 16942 2564 16948 2576
rect 16347 2536 16948 2564
rect 16347 2533 16359 2536
rect 16301 2527 16359 2533
rect 16942 2524 16948 2536
rect 17000 2524 17006 2576
rect 17865 2567 17923 2573
rect 17865 2533 17877 2567
rect 17911 2564 17923 2567
rect 18414 2564 18420 2576
rect 17911 2536 18420 2564
rect 17911 2533 17923 2536
rect 17865 2527 17923 2533
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18969 2567 19027 2573
rect 18969 2533 18981 2567
rect 19015 2564 19027 2567
rect 19610 2564 19616 2576
rect 19015 2536 19616 2564
rect 19015 2533 19027 2536
rect 18969 2527 19027 2533
rect 19610 2524 19616 2536
rect 19668 2524 19674 2576
rect 19720 2564 19748 2604
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 20622 2632 20628 2644
rect 20036 2604 20628 2632
rect 20036 2592 20042 2604
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 21266 2632 21272 2644
rect 20824 2604 21272 2632
rect 20162 2564 20168 2576
rect 19720 2536 20168 2564
rect 20162 2524 20168 2536
rect 20220 2524 20226 2576
rect 20824 2564 20852 2604
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 22002 2632 22008 2644
rect 21963 2604 22008 2632
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22112 2604 23336 2632
rect 20364 2536 20852 2564
rect 20892 2567 20950 2573
rect 1854 2496 1860 2508
rect 1815 2468 1860 2496
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 2832 2468 2881 2496
rect 2832 2456 2838 2468
rect 2869 2465 2881 2468
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4614 2496 4620 2508
rect 4387 2468 4620 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2496 5043 2499
rect 5074 2496 5080 2508
rect 5031 2468 5080 2496
rect 5031 2465 5043 2468
rect 4985 2459 5043 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 5994 2496 6000 2508
rect 5859 2468 6000 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6454 2456 6460 2508
rect 6512 2496 6518 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 6512 2468 7021 2496
rect 6512 2456 6518 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 8018 2496 8024 2508
rect 7791 2468 8024 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2496 8542 2508
rect 9582 2496 9588 2508
rect 8536 2468 9588 2496
rect 8536 2456 8542 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 11514 2496 11520 2508
rect 11195 2468 11520 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11514 2456 11520 2468
rect 11572 2456 11578 2508
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11940 2468 12265 2496
rect 11940 2456 11946 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 12483 2468 12572 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 11238 2428 11244 2440
rect 5184 2400 11244 2428
rect 5184 2369 5212 2400
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2428 11391 2431
rect 12544 2428 12572 2468
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 13814 2496 13820 2508
rect 12676 2468 12721 2496
rect 13775 2468 13820 2496
rect 12676 2456 12682 2468
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 14274 2456 14280 2508
rect 14332 2496 14338 2508
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 14332 2468 15025 2496
rect 14332 2456 14338 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 16022 2496 16028 2508
rect 15983 2468 16028 2496
rect 15013 2459 15071 2465
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16390 2496 16396 2508
rect 16351 2468 16396 2496
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 17494 2456 17500 2508
rect 17552 2496 17558 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17552 2468 17693 2496
rect 17552 2456 17558 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 18785 2499 18843 2505
rect 18785 2465 18797 2499
rect 18831 2465 18843 2499
rect 18785 2459 18843 2465
rect 19061 2499 19119 2505
rect 19061 2465 19073 2499
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 19153 2499 19211 2505
rect 19153 2465 19165 2499
rect 19199 2496 19211 2499
rect 20364 2496 20392 2536
rect 20892 2533 20904 2567
rect 20938 2564 20950 2567
rect 21174 2564 21180 2576
rect 20938 2536 21180 2564
rect 20938 2533 20950 2536
rect 20892 2527 20950 2533
rect 21174 2524 21180 2536
rect 21232 2524 21238 2576
rect 21284 2564 21312 2592
rect 22112 2564 22140 2604
rect 23198 2564 23204 2576
rect 21284 2536 22140 2564
rect 23159 2536 23204 2564
rect 23198 2524 23204 2536
rect 23256 2524 23262 2576
rect 19199 2468 20392 2496
rect 19199 2465 19211 2468
rect 19153 2459 19211 2465
rect 11379 2400 12434 2428
rect 12544 2400 15148 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 3053 2363 3111 2369
rect 3053 2329 3065 2363
rect 3099 2360 3111 2363
rect 5169 2363 5227 2369
rect 3099 2332 5120 2360
rect 3099 2329 3111 2332
rect 3053 2323 3111 2329
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 5092 2292 5120 2332
rect 5169 2329 5181 2363
rect 5215 2329 5227 2363
rect 7742 2360 7748 2372
rect 5169 2323 5227 2329
rect 5276 2332 7748 2360
rect 5276 2292 5304 2332
rect 7742 2320 7748 2332
rect 7800 2320 7806 2372
rect 7929 2363 7987 2369
rect 7929 2329 7941 2363
rect 7975 2360 7987 2363
rect 8294 2360 8300 2372
rect 7975 2332 8300 2360
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9674 2360 9680 2372
rect 8711 2332 9680 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 10594 2360 10600 2372
rect 10555 2332 10600 2360
rect 10594 2320 10600 2332
rect 10652 2320 10658 2372
rect 12406 2360 12434 2400
rect 15010 2360 15016 2372
rect 12406 2332 15016 2360
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 5092 2264 5304 2292
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 9766 2292 9772 2304
rect 7147 2264 9772 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 13906 2292 13912 2304
rect 13867 2264 13912 2292
rect 13906 2252 13912 2264
rect 13964 2252 13970 2304
rect 15120 2292 15148 2400
rect 15197 2363 15255 2369
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 17126 2360 17132 2372
rect 15243 2332 17132 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 18800 2360 18828 2459
rect 19076 2428 19104 2459
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 20625 2499 20683 2505
rect 20625 2496 20637 2499
rect 20496 2468 20637 2496
rect 20496 2456 20502 2468
rect 20625 2465 20637 2468
rect 20671 2465 20683 2499
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 20625 2459 20683 2465
rect 20732 2468 22937 2496
rect 19978 2428 19984 2440
rect 19076 2400 19984 2428
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20732 2428 20760 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 23106 2496 23112 2508
rect 23067 2468 23112 2496
rect 22925 2459 22983 2465
rect 23106 2456 23112 2468
rect 23164 2456 23170 2508
rect 23308 2505 23336 2604
rect 23382 2592 23388 2644
rect 23440 2632 23446 2644
rect 23477 2635 23535 2641
rect 23477 2632 23489 2635
rect 23440 2604 23489 2632
rect 23440 2592 23446 2604
rect 23477 2601 23489 2604
rect 23523 2601 23535 2635
rect 23477 2595 23535 2601
rect 24762 2592 24768 2644
rect 24820 2632 24826 2644
rect 25777 2635 25835 2641
rect 25777 2632 25789 2635
rect 24820 2604 25789 2632
rect 24820 2592 24826 2604
rect 25777 2601 25789 2604
rect 25823 2601 25835 2635
rect 25777 2595 25835 2601
rect 25866 2592 25872 2644
rect 25924 2632 25930 2644
rect 27249 2635 27307 2641
rect 27249 2632 27261 2635
rect 25924 2604 27261 2632
rect 25924 2592 25930 2604
rect 27249 2601 27261 2604
rect 27295 2601 27307 2635
rect 27249 2595 27307 2601
rect 24486 2524 24492 2576
rect 24544 2564 24550 2576
rect 25685 2567 25743 2573
rect 25685 2564 25697 2567
rect 24544 2536 25697 2564
rect 24544 2524 24550 2536
rect 25685 2533 25697 2536
rect 25731 2533 25743 2567
rect 25685 2527 25743 2533
rect 26421 2567 26479 2573
rect 26421 2533 26433 2567
rect 26467 2564 26479 2567
rect 27062 2564 27068 2576
rect 26467 2536 27068 2564
rect 26467 2533 26479 2536
rect 26421 2527 26479 2533
rect 27062 2524 27068 2536
rect 27120 2524 27126 2576
rect 23293 2499 23351 2505
rect 23293 2465 23305 2499
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 24029 2499 24087 2505
rect 24029 2465 24041 2499
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 27157 2499 27215 2505
rect 27157 2465 27169 2499
rect 27203 2496 27215 2499
rect 28534 2496 28540 2508
rect 27203 2468 28540 2496
rect 27203 2465 27215 2468
rect 27157 2459 27215 2465
rect 20548 2400 20760 2428
rect 20548 2372 20576 2400
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 24044 2428 24072 2459
rect 28534 2456 28540 2468
rect 28592 2456 28598 2508
rect 23072 2400 24072 2428
rect 23072 2388 23078 2400
rect 20530 2360 20536 2372
rect 18800 2332 20536 2360
rect 20530 2320 20536 2332
rect 20588 2320 20594 2372
rect 24946 2360 24952 2372
rect 22066 2332 24952 2360
rect 22066 2292 22094 2332
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 26605 2363 26663 2369
rect 26605 2329 26617 2363
rect 26651 2360 26663 2363
rect 28074 2360 28080 2372
rect 26651 2332 28080 2360
rect 26651 2329 26663 2332
rect 26605 2323 26663 2329
rect 28074 2320 28080 2332
rect 28132 2320 28138 2372
rect 24118 2292 24124 2304
rect 15120 2264 22094 2292
rect 24079 2264 24124 2292
rect 24118 2252 24124 2264
rect 24176 2252 24182 2304
rect 1104 2202 28428 2224
rect 1104 2150 5536 2202
rect 5588 2150 5600 2202
rect 5652 2150 5664 2202
rect 5716 2150 5728 2202
rect 5780 2150 14644 2202
rect 14696 2150 14708 2202
rect 14760 2150 14772 2202
rect 14824 2150 14836 2202
rect 14888 2150 23752 2202
rect 23804 2150 23816 2202
rect 23868 2150 23880 2202
rect 23932 2150 23944 2202
rect 23996 2150 28428 2202
rect 1104 2128 28428 2150
rect 11238 2048 11244 2100
rect 11296 2088 11302 2100
rect 17678 2088 17684 2100
rect 11296 2060 17684 2088
rect 11296 2048 11302 2060
rect 17678 2048 17684 2060
rect 17736 2048 17742 2100
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 23106 2020 23112 2032
rect 4120 1992 23112 2020
rect 4120 1980 4126 1992
rect 23106 1980 23112 1992
rect 23164 1980 23170 2032
rect 8202 1912 8208 1964
rect 8260 1952 8266 1964
rect 24118 1952 24124 1964
rect 8260 1924 24124 1952
rect 8260 1912 8266 1924
rect 24118 1912 24124 1924
rect 24176 1912 24182 1964
rect 1946 1844 1952 1896
rect 2004 1884 2010 1896
rect 10502 1884 10508 1896
rect 2004 1856 10508 1884
rect 2004 1844 2010 1856
rect 10502 1844 10508 1856
rect 10560 1844 10566 1896
rect 13906 1844 13912 1896
rect 13964 1884 13970 1896
rect 22186 1884 22192 1896
rect 13964 1856 22192 1884
rect 13964 1844 13970 1856
rect 22186 1844 22192 1856
rect 22244 1844 22250 1896
rect 7742 1776 7748 1828
rect 7800 1816 7806 1828
rect 7800 1788 12434 1816
rect 7800 1776 7806 1788
rect 12406 1748 12434 1788
rect 15010 1776 15016 1828
rect 15068 1816 15074 1828
rect 21910 1816 21916 1828
rect 15068 1788 21916 1816
rect 15068 1776 15074 1788
rect 21910 1776 21916 1788
rect 21968 1776 21974 1828
rect 18690 1748 18696 1760
rect 12406 1720 18696 1748
rect 18690 1708 18696 1720
rect 18748 1708 18754 1760
<< via1 >>
rect 15568 29656 15620 29708
rect 27344 29656 27396 29708
rect 9956 29520 10008 29572
rect 20076 29520 20128 29572
rect 15844 29452 15896 29504
rect 21272 29452 21324 29504
rect 5536 29350 5588 29402
rect 5600 29350 5652 29402
rect 5664 29350 5716 29402
rect 5728 29350 5780 29402
rect 14644 29350 14696 29402
rect 14708 29350 14760 29402
rect 14772 29350 14824 29402
rect 14836 29350 14888 29402
rect 23752 29350 23804 29402
rect 23816 29350 23868 29402
rect 23880 29350 23932 29402
rect 23944 29350 23996 29402
rect 3700 29248 3752 29300
rect 6000 29248 6052 29300
rect 7840 29291 7892 29300
rect 7840 29257 7849 29291
rect 7849 29257 7883 29291
rect 7883 29257 7892 29291
rect 7840 29248 7892 29257
rect 10600 29248 10652 29300
rect 12532 29248 12584 29300
rect 15752 29248 15804 29300
rect 17960 29248 18012 29300
rect 20720 29248 20772 29300
rect 21180 29248 21232 29300
rect 22100 29248 22152 29300
rect 28080 29248 28132 29300
rect 2412 29180 2464 29232
rect 5908 29180 5960 29232
rect 8760 29180 8812 29232
rect 18880 29180 18932 29232
rect 19800 29180 19852 29232
rect 27620 29180 27672 29232
rect 2964 29112 3016 29164
rect 1860 29087 1912 29096
rect 1860 29053 1869 29087
rect 1869 29053 1903 29087
rect 1903 29053 1912 29087
rect 1860 29044 1912 29053
rect 1952 29044 2004 29096
rect 9956 29087 10008 29096
rect 2228 28976 2280 29028
rect 5356 28976 5408 29028
rect 5632 29019 5684 29028
rect 5632 28985 5641 29019
rect 5641 28985 5675 29019
rect 5675 28985 5684 29019
rect 5632 28976 5684 28985
rect 7748 29019 7800 29028
rect 7748 28985 7757 29019
rect 7757 28985 7791 29019
rect 7791 28985 7800 29019
rect 7748 28976 7800 28985
rect 9956 29053 9965 29087
rect 9965 29053 9999 29087
rect 9999 29053 10008 29087
rect 9956 29044 10008 29053
rect 10968 29044 11020 29096
rect 12440 29044 12492 29096
rect 12900 29044 12952 29096
rect 15016 29087 15068 29096
rect 15016 29053 15025 29087
rect 15025 29053 15059 29087
rect 15059 29053 15068 29087
rect 15016 29044 15068 29053
rect 16304 29044 16356 29096
rect 17040 29044 17092 29096
rect 17684 29044 17736 29096
rect 18052 29044 18104 29096
rect 19708 29112 19760 29164
rect 27344 29155 27396 29164
rect 6920 28908 6972 28960
rect 8300 28908 8352 28960
rect 9864 28976 9916 29028
rect 10692 29019 10744 29028
rect 9496 28908 9548 28960
rect 10692 28985 10701 29019
rect 10701 28985 10735 29019
rect 10735 28985 10744 29019
rect 10692 28976 10744 28985
rect 12808 28976 12860 29028
rect 15844 28976 15896 29028
rect 16028 28908 16080 28960
rect 18788 28976 18840 29028
rect 21640 29044 21692 29096
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 25964 29044 26016 29096
rect 26148 29044 26200 29096
rect 27160 29087 27212 29096
rect 27160 29053 27169 29087
rect 27169 29053 27203 29087
rect 27203 29053 27212 29087
rect 27160 29044 27212 29053
rect 23756 29019 23808 29028
rect 18144 28951 18196 28960
rect 18144 28917 18153 28951
rect 18153 28917 18187 28951
rect 18187 28917 18196 28951
rect 18144 28908 18196 28917
rect 20996 28908 21048 28960
rect 23756 28985 23765 29019
rect 23765 28985 23799 29019
rect 23799 28985 23808 29019
rect 23756 28976 23808 28985
rect 25596 28976 25648 29028
rect 26792 28976 26844 29028
rect 24584 28908 24636 28960
rect 10090 28806 10142 28858
rect 10154 28806 10206 28858
rect 10218 28806 10270 28858
rect 10282 28806 10334 28858
rect 19198 28806 19250 28858
rect 19262 28806 19314 28858
rect 19326 28806 19378 28858
rect 19390 28806 19442 28858
rect 480 28704 532 28756
rect 2320 28704 2372 28756
rect 5632 28704 5684 28756
rect 1768 28568 1820 28620
rect 3424 28568 3476 28620
rect 4160 28568 4212 28620
rect 5080 28611 5132 28620
rect 5080 28577 5089 28611
rect 5089 28577 5123 28611
rect 5123 28577 5132 28611
rect 5080 28568 5132 28577
rect 7472 28679 7524 28688
rect 7472 28645 7481 28679
rect 7481 28645 7515 28679
rect 7515 28645 7524 28679
rect 7472 28636 7524 28645
rect 9680 28636 9732 28688
rect 7104 28568 7156 28620
rect 7564 28611 7616 28620
rect 7564 28577 7573 28611
rect 7573 28577 7607 28611
rect 7607 28577 7616 28611
rect 7564 28568 7616 28577
rect 7840 28568 7892 28620
rect 8300 28611 8352 28620
rect 8300 28577 8309 28611
rect 8309 28577 8343 28611
rect 8343 28577 8352 28611
rect 8300 28568 8352 28577
rect 9496 28611 9548 28620
rect 9496 28577 9505 28611
rect 9505 28577 9539 28611
rect 9539 28577 9548 28611
rect 9496 28568 9548 28577
rect 10508 28611 10560 28620
rect 10508 28577 10542 28611
rect 10542 28577 10560 28611
rect 11060 28636 11112 28688
rect 16028 28704 16080 28756
rect 16396 28704 16448 28756
rect 10508 28568 10560 28577
rect 17592 28636 17644 28688
rect 20260 28636 20312 28688
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 16028 28568 16080 28620
rect 16120 28568 16172 28620
rect 18052 28568 18104 28620
rect 20076 28611 20128 28620
rect 20076 28577 20085 28611
rect 20085 28577 20119 28611
rect 20119 28577 20128 28611
rect 20076 28568 20128 28577
rect 20996 28568 21048 28620
rect 24400 28636 24452 28688
rect 29000 28636 29052 28688
rect 8576 28500 8628 28552
rect 9956 28500 10008 28552
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 14464 28500 14516 28552
rect 17224 28500 17276 28552
rect 20904 28500 20956 28552
rect 23480 28568 23532 28620
rect 24216 28568 24268 28620
rect 25044 28568 25096 28620
rect 23756 28500 23808 28552
rect 26424 28568 26476 28620
rect 9864 28432 9916 28484
rect 4988 28364 5040 28416
rect 7472 28364 7524 28416
rect 10416 28364 10468 28416
rect 11152 28364 11204 28416
rect 17408 28432 17460 28484
rect 17500 28364 17552 28416
rect 18880 28407 18932 28416
rect 18880 28373 18889 28407
rect 18889 28373 18923 28407
rect 18923 28373 18932 28407
rect 18880 28364 18932 28373
rect 22652 28364 22704 28416
rect 26148 28364 26200 28416
rect 5536 28262 5588 28314
rect 5600 28262 5652 28314
rect 5664 28262 5716 28314
rect 5728 28262 5780 28314
rect 14644 28262 14696 28314
rect 14708 28262 14760 28314
rect 14772 28262 14824 28314
rect 14836 28262 14888 28314
rect 23752 28262 23804 28314
rect 23816 28262 23868 28314
rect 23880 28262 23932 28314
rect 23944 28262 23996 28314
rect 2780 28092 2832 28144
rect 2964 28135 3016 28144
rect 2964 28101 2973 28135
rect 2973 28101 3007 28135
rect 3007 28101 3016 28135
rect 2964 28092 3016 28101
rect 10416 28092 10468 28144
rect 12992 28092 13044 28144
rect 18788 28092 18840 28144
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 2136 27999 2188 28008
rect 2136 27965 2145 27999
rect 2145 27965 2179 27999
rect 2179 27965 2188 27999
rect 2136 27956 2188 27965
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 2780 27956 2832 27965
rect 7472 27956 7524 28008
rect 9496 27956 9548 28008
rect 10232 28024 10284 28076
rect 8760 27888 8812 27940
rect 9680 27888 9732 27940
rect 10692 27956 10744 28008
rect 11520 27956 11572 28008
rect 14372 27999 14424 28008
rect 14372 27965 14381 27999
rect 14381 27965 14415 27999
rect 14415 27965 14424 27999
rect 14372 27956 14424 27965
rect 15200 27956 15252 28008
rect 17224 27956 17276 28008
rect 18144 27956 18196 28008
rect 19708 27956 19760 28008
rect 21732 28024 21784 28076
rect 21272 27999 21324 28008
rect 15292 27888 15344 27940
rect 17684 27888 17736 27940
rect 4436 27820 4488 27872
rect 6644 27820 6696 27872
rect 7564 27820 7616 27872
rect 9772 27820 9824 27872
rect 10416 27820 10468 27872
rect 13084 27820 13136 27872
rect 15384 27820 15436 27872
rect 16120 27820 16172 27872
rect 17960 27820 18012 27872
rect 21272 27965 21281 27999
rect 21281 27965 21315 27999
rect 21315 27965 21324 27999
rect 21272 27956 21324 27965
rect 21640 27956 21692 28008
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 24124 27956 24176 28008
rect 24584 27999 24636 28008
rect 24584 27965 24593 27999
rect 24593 27965 24627 27999
rect 24627 27965 24636 27999
rect 24584 27956 24636 27965
rect 25320 27999 25372 28008
rect 25320 27965 25329 27999
rect 25329 27965 25363 27999
rect 25363 27965 25372 27999
rect 25320 27956 25372 27965
rect 25964 27999 26016 28008
rect 25964 27965 25973 27999
rect 25973 27965 26007 27999
rect 26007 27965 26016 27999
rect 25964 27956 26016 27965
rect 26240 27956 26292 28008
rect 20812 27863 20864 27872
rect 20812 27829 20821 27863
rect 20821 27829 20855 27863
rect 20855 27829 20864 27863
rect 20812 27820 20864 27829
rect 22376 27820 22428 27872
rect 24676 27820 24728 27872
rect 10090 27718 10142 27770
rect 10154 27718 10206 27770
rect 10218 27718 10270 27770
rect 10282 27718 10334 27770
rect 19198 27718 19250 27770
rect 19262 27718 19314 27770
rect 19326 27718 19378 27770
rect 19390 27718 19442 27770
rect 10508 27616 10560 27668
rect 940 27548 992 27600
rect 2780 27548 2832 27600
rect 7380 27548 7432 27600
rect 2872 27480 2924 27532
rect 7656 27480 7708 27532
rect 9864 27548 9916 27600
rect 12256 27616 12308 27668
rect 10968 27548 11020 27600
rect 14280 27548 14332 27600
rect 9772 27480 9824 27532
rect 5172 27412 5224 27464
rect 9404 27412 9456 27464
rect 10508 27523 10560 27532
rect 10508 27489 10517 27523
rect 10517 27489 10551 27523
rect 10551 27489 10560 27523
rect 10508 27480 10560 27489
rect 12624 27480 12676 27532
rect 13360 27480 13412 27532
rect 15108 27616 15160 27668
rect 15292 27659 15344 27668
rect 15292 27625 15301 27659
rect 15301 27625 15335 27659
rect 15335 27625 15344 27659
rect 15292 27616 15344 27625
rect 16028 27616 16080 27668
rect 18052 27659 18104 27668
rect 18052 27625 18061 27659
rect 18061 27625 18095 27659
rect 18095 27625 18104 27659
rect 18052 27616 18104 27625
rect 15384 27548 15436 27600
rect 15568 27548 15620 27600
rect 15108 27523 15160 27532
rect 11060 27412 11112 27464
rect 11888 27455 11940 27464
rect 11888 27421 11897 27455
rect 11897 27421 11931 27455
rect 11931 27421 11940 27455
rect 11888 27412 11940 27421
rect 14372 27412 14424 27464
rect 15108 27489 15117 27523
rect 15117 27489 15151 27523
rect 15151 27489 15160 27523
rect 15108 27480 15160 27489
rect 15200 27480 15252 27532
rect 15844 27480 15896 27532
rect 16396 27548 16448 27600
rect 17408 27548 17460 27600
rect 18328 27548 18380 27600
rect 18880 27548 18932 27600
rect 20812 27548 20864 27600
rect 25780 27591 25832 27600
rect 25780 27557 25789 27591
rect 25789 27557 25823 27591
rect 25823 27557 25832 27591
rect 25780 27548 25832 27557
rect 26056 27548 26108 27600
rect 16580 27480 16632 27532
rect 17960 27480 18012 27532
rect 18420 27480 18472 27532
rect 24308 27480 24360 27532
rect 7564 27344 7616 27396
rect 17684 27412 17736 27464
rect 20352 27455 20404 27464
rect 20352 27421 20361 27455
rect 20361 27421 20395 27455
rect 20395 27421 20404 27455
rect 20352 27412 20404 27421
rect 26424 27480 26476 27532
rect 27344 27480 27396 27532
rect 26516 27412 26568 27464
rect 2964 27276 3016 27328
rect 7380 27276 7432 27328
rect 8668 27276 8720 27328
rect 17500 27344 17552 27396
rect 21732 27387 21784 27396
rect 21732 27353 21741 27387
rect 21741 27353 21775 27387
rect 21775 27353 21784 27387
rect 21732 27344 21784 27353
rect 13084 27276 13136 27328
rect 13268 27319 13320 27328
rect 13268 27285 13277 27319
rect 13277 27285 13311 27319
rect 13311 27285 13320 27319
rect 13268 27276 13320 27285
rect 16948 27319 17000 27328
rect 16948 27285 16957 27319
rect 16957 27285 16991 27319
rect 16991 27285 17000 27319
rect 16948 27276 17000 27285
rect 18696 27319 18748 27328
rect 18696 27285 18705 27319
rect 18705 27285 18739 27319
rect 18739 27285 18748 27319
rect 18696 27276 18748 27285
rect 5536 27174 5588 27226
rect 5600 27174 5652 27226
rect 5664 27174 5716 27226
rect 5728 27174 5780 27226
rect 14644 27174 14696 27226
rect 14708 27174 14760 27226
rect 14772 27174 14824 27226
rect 14836 27174 14888 27226
rect 23752 27174 23804 27226
rect 23816 27174 23868 27226
rect 23880 27174 23932 27226
rect 23944 27174 23996 27226
rect 7656 27115 7708 27124
rect 7656 27081 7665 27115
rect 7665 27081 7699 27115
rect 7699 27081 7708 27115
rect 7656 27072 7708 27081
rect 8760 27072 8812 27124
rect 18696 27072 18748 27124
rect 2136 26911 2188 26920
rect 2136 26877 2145 26911
rect 2145 26877 2179 26911
rect 2179 26877 2188 26911
rect 2136 26868 2188 26877
rect 7104 26911 7156 26920
rect 7104 26877 7113 26911
rect 7113 26877 7147 26911
rect 7147 26877 7156 26911
rect 7104 26868 7156 26877
rect 7380 26911 7432 26920
rect 7380 26877 7389 26911
rect 7389 26877 7423 26911
rect 7423 26877 7432 26911
rect 7380 26868 7432 26877
rect 7840 26868 7892 26920
rect 9220 26936 9272 26988
rect 9864 27004 9916 27056
rect 10048 27004 10100 27056
rect 7564 26800 7616 26852
rect 9404 26868 9456 26920
rect 9680 26800 9732 26852
rect 9588 26732 9640 26784
rect 10140 26868 10192 26920
rect 11888 26868 11940 26920
rect 13360 26868 13412 26920
rect 10508 26800 10560 26852
rect 12716 26800 12768 26852
rect 9860 26732 9912 26784
rect 9956 26732 10008 26784
rect 12532 26732 12584 26784
rect 15108 26868 15160 26920
rect 15568 26936 15620 26988
rect 16028 26936 16080 26988
rect 15476 26868 15528 26920
rect 16396 27004 16448 27056
rect 26884 27047 26936 27056
rect 26884 27013 26893 27047
rect 26893 27013 26927 27047
rect 26927 27013 26936 27047
rect 26884 27004 26936 27013
rect 16212 26936 16264 26988
rect 16396 26868 16448 26920
rect 17500 26911 17552 26920
rect 17500 26877 17509 26911
rect 17509 26877 17543 26911
rect 17543 26877 17552 26911
rect 17500 26868 17552 26877
rect 18328 26911 18380 26920
rect 18328 26877 18337 26911
rect 18337 26877 18371 26911
rect 18371 26877 18380 26911
rect 18328 26868 18380 26877
rect 18788 26868 18840 26920
rect 21732 26868 21784 26920
rect 21824 26868 21876 26920
rect 22928 26868 22980 26920
rect 24308 26868 24360 26920
rect 16672 26800 16724 26852
rect 18236 26800 18288 26852
rect 14188 26732 14240 26784
rect 15568 26775 15620 26784
rect 15568 26741 15577 26775
rect 15577 26741 15611 26775
rect 15611 26741 15620 26775
rect 15568 26732 15620 26741
rect 16580 26732 16632 26784
rect 17868 26775 17920 26784
rect 17868 26741 17877 26775
rect 17877 26741 17911 26775
rect 17911 26741 17920 26775
rect 17868 26732 17920 26741
rect 18512 26732 18564 26784
rect 18604 26732 18656 26784
rect 21548 26775 21600 26784
rect 21548 26741 21557 26775
rect 21557 26741 21591 26775
rect 21591 26741 21600 26775
rect 21548 26732 21600 26741
rect 23296 26800 23348 26852
rect 23204 26732 23256 26784
rect 23388 26775 23440 26784
rect 23388 26741 23397 26775
rect 23397 26741 23431 26775
rect 23431 26741 23440 26775
rect 23388 26732 23440 26741
rect 10090 26630 10142 26682
rect 10154 26630 10206 26682
rect 10218 26630 10270 26682
rect 10282 26630 10334 26682
rect 19198 26630 19250 26682
rect 19262 26630 19314 26682
rect 19326 26630 19378 26682
rect 19390 26630 19442 26682
rect 1952 26571 2004 26580
rect 1952 26537 1961 26571
rect 1961 26537 1995 26571
rect 1995 26537 2004 26571
rect 1952 26528 2004 26537
rect 9496 26528 9548 26580
rect 9956 26460 10008 26512
rect 16672 26528 16724 26580
rect 18236 26528 18288 26580
rect 18788 26528 18840 26580
rect 22284 26571 22336 26580
rect 22284 26537 22293 26571
rect 22293 26537 22327 26571
rect 22327 26537 22336 26571
rect 22284 26528 22336 26537
rect 23296 26528 23348 26580
rect 24308 26571 24360 26580
rect 24308 26537 24317 26571
rect 24317 26537 24351 26571
rect 24351 26537 24360 26571
rect 24308 26528 24360 26537
rect 2136 26392 2188 26444
rect 11060 26392 11112 26444
rect 11888 26460 11940 26512
rect 13728 26460 13780 26512
rect 15568 26460 15620 26512
rect 17868 26460 17920 26512
rect 23388 26460 23440 26512
rect 27436 26460 27488 26512
rect 27712 26503 27764 26512
rect 27712 26469 27721 26503
rect 27721 26469 27755 26503
rect 27755 26469 27764 26503
rect 27712 26460 27764 26469
rect 9496 26367 9548 26376
rect 9496 26333 9505 26367
rect 9505 26333 9539 26367
rect 9539 26333 9548 26367
rect 9496 26324 9548 26333
rect 2136 26188 2188 26240
rect 9864 26188 9916 26240
rect 12164 26188 12216 26240
rect 13268 26392 13320 26444
rect 14464 26392 14516 26444
rect 17224 26392 17276 26444
rect 20352 26392 20404 26444
rect 21456 26392 21508 26444
rect 27160 26392 27212 26444
rect 22836 26324 22888 26376
rect 14464 26256 14516 26308
rect 26976 26299 27028 26308
rect 26976 26265 26985 26299
rect 26985 26265 27019 26299
rect 27019 26265 27028 26299
rect 26976 26256 27028 26265
rect 13176 26231 13228 26240
rect 13176 26197 13185 26231
rect 13185 26197 13219 26231
rect 13219 26197 13228 26231
rect 13176 26188 13228 26197
rect 5536 26086 5588 26138
rect 5600 26086 5652 26138
rect 5664 26086 5716 26138
rect 5728 26086 5780 26138
rect 14644 26086 14696 26138
rect 14708 26086 14760 26138
rect 14772 26086 14824 26138
rect 14836 26086 14888 26138
rect 23752 26086 23804 26138
rect 23816 26086 23868 26138
rect 23880 26086 23932 26138
rect 23944 26086 23996 26138
rect 12348 25984 12400 26036
rect 12624 26027 12676 26036
rect 12624 25993 12633 26027
rect 12633 25993 12667 26027
rect 12667 25993 12676 26027
rect 12624 25984 12676 25993
rect 21456 26027 21508 26036
rect 8208 25916 8260 25968
rect 14280 25916 14332 25968
rect 1676 25891 1728 25900
rect 1676 25857 1685 25891
rect 1685 25857 1719 25891
rect 1719 25857 1728 25891
rect 1676 25848 1728 25857
rect 2136 25823 2188 25832
rect 2136 25789 2145 25823
rect 2145 25789 2179 25823
rect 2179 25789 2188 25823
rect 2136 25780 2188 25789
rect 2872 25823 2924 25832
rect 2872 25789 2881 25823
rect 2881 25789 2915 25823
rect 2915 25789 2924 25823
rect 2872 25780 2924 25789
rect 5264 25823 5316 25832
rect 5264 25789 5273 25823
rect 5273 25789 5307 25823
rect 5307 25789 5316 25823
rect 5264 25780 5316 25789
rect 5908 25780 5960 25832
rect 7380 25780 7432 25832
rect 7472 25780 7524 25832
rect 9496 25780 9548 25832
rect 11244 25848 11296 25900
rect 14464 25891 14516 25900
rect 10416 25780 10468 25832
rect 12072 25823 12124 25832
rect 12072 25789 12081 25823
rect 12081 25789 12115 25823
rect 12115 25789 12124 25823
rect 12072 25780 12124 25789
rect 12164 25780 12216 25832
rect 3332 25712 3384 25764
rect 11428 25712 11480 25764
rect 12256 25755 12308 25764
rect 12256 25721 12265 25755
rect 12265 25721 12299 25755
rect 12299 25721 12308 25755
rect 13636 25780 13688 25832
rect 14096 25780 14148 25832
rect 12256 25712 12308 25721
rect 14004 25712 14056 25764
rect 14464 25857 14473 25891
rect 14473 25857 14507 25891
rect 14507 25857 14516 25891
rect 14464 25848 14516 25857
rect 16396 25916 16448 25968
rect 21456 25993 21465 26027
rect 21465 25993 21499 26027
rect 21499 25993 21508 26027
rect 21456 25984 21508 25993
rect 24216 26027 24268 26036
rect 24216 25993 24225 26027
rect 24225 25993 24259 26027
rect 24259 25993 24268 26027
rect 24216 25984 24268 25993
rect 26884 25891 26936 25900
rect 15660 25780 15712 25832
rect 16028 25823 16080 25832
rect 16028 25789 16037 25823
rect 16037 25789 16071 25823
rect 16071 25789 16080 25823
rect 16028 25780 16080 25789
rect 16212 25823 16264 25832
rect 16212 25789 16221 25823
rect 16221 25789 16255 25823
rect 16255 25789 16264 25823
rect 16212 25780 16264 25789
rect 17224 25780 17276 25832
rect 20904 25823 20956 25832
rect 4252 25687 4304 25696
rect 4252 25653 4261 25687
rect 4261 25653 4295 25687
rect 4295 25653 4304 25687
rect 4252 25644 4304 25653
rect 5816 25687 5868 25696
rect 5816 25653 5825 25687
rect 5825 25653 5859 25687
rect 5859 25653 5868 25687
rect 5816 25644 5868 25653
rect 6092 25644 6144 25696
rect 11152 25687 11204 25696
rect 11152 25653 11161 25687
rect 11161 25653 11195 25687
rect 11195 25653 11204 25687
rect 11152 25644 11204 25653
rect 12624 25644 12676 25696
rect 14280 25644 14332 25696
rect 16028 25644 16080 25696
rect 20904 25789 20913 25823
rect 20913 25789 20947 25823
rect 20947 25789 20956 25823
rect 20904 25780 20956 25789
rect 22284 25780 22336 25832
rect 22836 25823 22888 25832
rect 22836 25789 22845 25823
rect 22845 25789 22879 25823
rect 22879 25789 22888 25823
rect 22836 25780 22888 25789
rect 26884 25857 26893 25891
rect 26893 25857 26927 25891
rect 26927 25857 26936 25891
rect 26884 25848 26936 25857
rect 26608 25780 26660 25832
rect 21088 25755 21140 25764
rect 21088 25721 21097 25755
rect 21097 25721 21131 25755
rect 21131 25721 21140 25755
rect 21088 25712 21140 25721
rect 18880 25644 18932 25696
rect 22284 25644 22336 25696
rect 22928 25644 22980 25696
rect 23388 25712 23440 25764
rect 24768 25712 24820 25764
rect 24952 25755 25004 25764
rect 24952 25721 24961 25755
rect 24961 25721 24995 25755
rect 24995 25721 25004 25755
rect 24952 25712 25004 25721
rect 24124 25644 24176 25696
rect 25228 25687 25280 25696
rect 25228 25653 25237 25687
rect 25237 25653 25271 25687
rect 25271 25653 25280 25687
rect 25228 25644 25280 25653
rect 10090 25542 10142 25594
rect 10154 25542 10206 25594
rect 10218 25542 10270 25594
rect 10282 25542 10334 25594
rect 19198 25542 19250 25594
rect 19262 25542 19314 25594
rect 19326 25542 19378 25594
rect 19390 25542 19442 25594
rect 3332 25483 3384 25492
rect 3332 25449 3341 25483
rect 3341 25449 3375 25483
rect 3375 25449 3384 25483
rect 3332 25440 3384 25449
rect 4252 25440 4304 25492
rect 2964 25415 3016 25424
rect 2964 25381 2973 25415
rect 2973 25381 3007 25415
rect 3007 25381 3016 25415
rect 2964 25372 3016 25381
rect 5816 25372 5868 25424
rect 7472 25440 7524 25492
rect 9680 25440 9732 25492
rect 10876 25440 10928 25492
rect 11428 25483 11480 25492
rect 11428 25449 11437 25483
rect 11437 25449 11471 25483
rect 11471 25449 11480 25483
rect 11428 25440 11480 25449
rect 12256 25440 12308 25492
rect 12716 25440 12768 25492
rect 13084 25440 13136 25492
rect 11152 25415 11204 25424
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 3148 25347 3200 25356
rect 2688 25236 2740 25288
rect 3148 25313 3157 25347
rect 3157 25313 3191 25347
rect 3191 25313 3200 25347
rect 3148 25304 3200 25313
rect 3332 25304 3384 25356
rect 5264 25304 5316 25356
rect 7104 25347 7156 25356
rect 7104 25313 7113 25347
rect 7113 25313 7147 25347
rect 7147 25313 7156 25347
rect 7104 25304 7156 25313
rect 7380 25347 7432 25356
rect 5172 25279 5224 25288
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 5172 25236 5224 25245
rect 7380 25313 7389 25347
rect 7389 25313 7423 25347
rect 7423 25313 7432 25347
rect 7380 25304 7432 25313
rect 7840 25304 7892 25356
rect 11152 25381 11161 25415
rect 11161 25381 11195 25415
rect 11195 25381 11204 25415
rect 11152 25372 11204 25381
rect 12532 25415 12584 25424
rect 12532 25381 12541 25415
rect 12541 25381 12575 25415
rect 12575 25381 12584 25415
rect 12532 25372 12584 25381
rect 13176 25372 13228 25424
rect 13728 25440 13780 25492
rect 13912 25440 13964 25492
rect 20904 25440 20956 25492
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 26608 25483 26660 25492
rect 26608 25449 26617 25483
rect 26617 25449 26651 25483
rect 26651 25449 26660 25483
rect 26608 25440 26660 25449
rect 9864 25304 9916 25356
rect 8024 25236 8076 25288
rect 10968 25304 11020 25356
rect 11244 25347 11296 25356
rect 11244 25313 11253 25347
rect 11253 25313 11287 25347
rect 11287 25313 11296 25347
rect 11244 25304 11296 25313
rect 12256 25347 12308 25356
rect 12256 25313 12265 25347
rect 12265 25313 12299 25347
rect 12299 25313 12308 25347
rect 12256 25304 12308 25313
rect 12808 25304 12860 25356
rect 13452 25347 13504 25356
rect 12072 25236 12124 25288
rect 10048 25168 10100 25220
rect 11888 25168 11940 25220
rect 12716 25236 12768 25288
rect 13084 25236 13136 25288
rect 13452 25313 13461 25347
rect 13461 25313 13495 25347
rect 13495 25313 13504 25347
rect 13452 25304 13504 25313
rect 13728 25304 13780 25356
rect 15200 25372 15252 25424
rect 23296 25372 23348 25424
rect 24952 25372 25004 25424
rect 25228 25372 25280 25424
rect 16672 25347 16724 25356
rect 16672 25313 16681 25347
rect 16681 25313 16715 25347
rect 16715 25313 16724 25347
rect 16672 25304 16724 25313
rect 17316 25347 17368 25356
rect 17316 25313 17325 25347
rect 17325 25313 17359 25347
rect 17359 25313 17368 25347
rect 17316 25304 17368 25313
rect 18144 25347 18196 25356
rect 13360 25236 13412 25288
rect 2136 25100 2188 25152
rect 4344 25143 4396 25152
rect 4344 25109 4353 25143
rect 4353 25109 4387 25143
rect 4387 25109 4396 25143
rect 4344 25100 4396 25109
rect 7656 25143 7708 25152
rect 7656 25109 7665 25143
rect 7665 25109 7699 25143
rect 7699 25109 7708 25143
rect 7656 25100 7708 25109
rect 8208 25143 8260 25152
rect 8208 25109 8217 25143
rect 8217 25109 8251 25143
rect 8251 25109 8260 25143
rect 8208 25100 8260 25109
rect 10140 25100 10192 25152
rect 10600 25100 10652 25152
rect 12256 25100 12308 25152
rect 12808 25100 12860 25152
rect 13728 25100 13780 25152
rect 17040 25168 17092 25220
rect 18144 25313 18153 25347
rect 18153 25313 18187 25347
rect 18187 25313 18196 25347
rect 18144 25304 18196 25313
rect 18788 25347 18840 25356
rect 18788 25313 18797 25347
rect 18797 25313 18831 25347
rect 18831 25313 18840 25347
rect 18788 25304 18840 25313
rect 22192 25304 22244 25356
rect 18696 25236 18748 25288
rect 24216 25304 24268 25356
rect 24768 25236 24820 25288
rect 26056 25304 26108 25356
rect 27160 25304 27212 25356
rect 21824 25168 21876 25220
rect 15108 25100 15160 25152
rect 16120 25143 16172 25152
rect 16120 25109 16129 25143
rect 16129 25109 16163 25143
rect 16163 25109 16172 25143
rect 16120 25100 16172 25109
rect 18328 25100 18380 25152
rect 5536 24998 5588 25050
rect 5600 24998 5652 25050
rect 5664 24998 5716 25050
rect 5728 24998 5780 25050
rect 14644 24998 14696 25050
rect 14708 24998 14760 25050
rect 14772 24998 14824 25050
rect 14836 24998 14888 25050
rect 23752 24998 23804 25050
rect 23816 24998 23868 25050
rect 23880 24998 23932 25050
rect 23944 24998 23996 25050
rect 4344 24896 4396 24948
rect 5264 24828 5316 24880
rect 7104 24828 7156 24880
rect 11428 24828 11480 24880
rect 12072 24828 12124 24880
rect 12624 24828 12676 24880
rect 13912 24828 13964 24880
rect 1492 24692 1544 24744
rect 2504 24760 2556 24812
rect 2688 24760 2740 24812
rect 2872 24760 2924 24812
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 3148 24692 3200 24744
rect 5172 24760 5224 24812
rect 10692 24760 10744 24812
rect 10048 24735 10100 24744
rect 3332 24624 3384 24676
rect 4804 24624 4856 24676
rect 1676 24599 1728 24608
rect 1676 24565 1685 24599
rect 1685 24565 1719 24599
rect 1719 24565 1728 24599
rect 1676 24556 1728 24565
rect 2780 24599 2832 24608
rect 2780 24565 2789 24599
rect 2789 24565 2823 24599
rect 2823 24565 2832 24599
rect 2780 24556 2832 24565
rect 4528 24556 4580 24608
rect 8576 24624 8628 24676
rect 8116 24556 8168 24608
rect 8944 24556 8996 24608
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 10140 24692 10192 24744
rect 10600 24735 10652 24744
rect 10600 24701 10609 24735
rect 10609 24701 10643 24735
rect 10643 24701 10652 24735
rect 10600 24692 10652 24701
rect 11060 24692 11112 24744
rect 13636 24760 13688 24812
rect 14004 24803 14056 24812
rect 14004 24769 14013 24803
rect 14013 24769 14047 24803
rect 14047 24769 14056 24803
rect 14004 24760 14056 24769
rect 14924 24828 14976 24880
rect 13084 24692 13136 24744
rect 13268 24735 13320 24744
rect 13268 24701 13277 24735
rect 13277 24701 13311 24735
rect 13311 24701 13320 24735
rect 13268 24692 13320 24701
rect 14188 24735 14240 24744
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 14280 24735 14332 24744
rect 14280 24701 14289 24735
rect 14289 24701 14323 24735
rect 14323 24701 14332 24735
rect 14280 24692 14332 24701
rect 15292 24735 15344 24744
rect 15292 24701 15301 24735
rect 15301 24701 15335 24735
rect 15335 24701 15344 24735
rect 15292 24692 15344 24701
rect 15660 24896 15712 24948
rect 18696 24896 18748 24948
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 19064 24828 19116 24880
rect 22100 24828 22152 24880
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 16212 24735 16264 24744
rect 16212 24701 16221 24735
rect 16221 24701 16255 24735
rect 16255 24701 16264 24735
rect 16212 24692 16264 24701
rect 10784 24624 10836 24676
rect 13544 24667 13596 24676
rect 13544 24633 13553 24667
rect 13553 24633 13587 24667
rect 13587 24633 13596 24667
rect 13544 24624 13596 24633
rect 17408 24692 17460 24744
rect 18144 24735 18196 24744
rect 18144 24701 18153 24735
rect 18153 24701 18187 24735
rect 18187 24701 18196 24735
rect 18144 24692 18196 24701
rect 18328 24735 18380 24744
rect 18328 24701 18337 24735
rect 18337 24701 18371 24735
rect 18371 24701 18380 24735
rect 18328 24692 18380 24701
rect 18880 24692 18932 24744
rect 21456 24692 21508 24744
rect 23204 24735 23256 24744
rect 23204 24701 23213 24735
rect 23213 24701 23247 24735
rect 23247 24701 23256 24735
rect 23204 24692 23256 24701
rect 23388 24735 23440 24744
rect 23388 24701 23397 24735
rect 23397 24701 23431 24735
rect 23431 24701 23440 24735
rect 23388 24692 23440 24701
rect 18972 24624 19024 24676
rect 21088 24624 21140 24676
rect 23296 24667 23348 24676
rect 23296 24633 23305 24667
rect 23305 24633 23339 24667
rect 23339 24633 23348 24667
rect 24124 24692 24176 24744
rect 26148 24735 26200 24744
rect 26148 24701 26157 24735
rect 26157 24701 26191 24735
rect 26191 24701 26200 24735
rect 26148 24692 26200 24701
rect 26608 24692 26660 24744
rect 23296 24624 23348 24633
rect 26332 24667 26384 24676
rect 26332 24633 26341 24667
rect 26341 24633 26375 24667
rect 26375 24633 26384 24667
rect 26332 24624 26384 24633
rect 26424 24667 26476 24676
rect 26424 24633 26433 24667
rect 26433 24633 26467 24667
rect 26467 24633 26476 24667
rect 26424 24624 26476 24633
rect 17500 24556 17552 24608
rect 22928 24556 22980 24608
rect 23388 24556 23440 24608
rect 26240 24556 26292 24608
rect 26700 24599 26752 24608
rect 26700 24565 26709 24599
rect 26709 24565 26743 24599
rect 26743 24565 26752 24599
rect 26700 24556 26752 24565
rect 10090 24454 10142 24506
rect 10154 24454 10206 24506
rect 10218 24454 10270 24506
rect 10282 24454 10334 24506
rect 19198 24454 19250 24506
rect 19262 24454 19314 24506
rect 19326 24454 19378 24506
rect 19390 24454 19442 24506
rect 3332 24395 3384 24404
rect 3332 24361 3341 24395
rect 3341 24361 3375 24395
rect 3375 24361 3384 24395
rect 3332 24352 3384 24361
rect 4804 24395 4856 24404
rect 2780 24284 2832 24336
rect 2872 24284 2924 24336
rect 3148 24284 3200 24336
rect 4528 24327 4580 24336
rect 4528 24293 4537 24327
rect 4537 24293 4571 24327
rect 4571 24293 4580 24327
rect 4528 24284 4580 24293
rect 4804 24361 4813 24395
rect 4813 24361 4847 24395
rect 4847 24361 4856 24395
rect 4804 24352 4856 24361
rect 4436 24259 4488 24268
rect 4436 24225 4445 24259
rect 4445 24225 4479 24259
rect 4479 24225 4488 24259
rect 4436 24216 4488 24225
rect 5908 24284 5960 24336
rect 7564 24352 7616 24404
rect 8576 24395 8628 24404
rect 8576 24361 8585 24395
rect 8585 24361 8619 24395
rect 8619 24361 8628 24395
rect 8576 24352 8628 24361
rect 13544 24352 13596 24404
rect 15200 24352 15252 24404
rect 15936 24352 15988 24404
rect 22652 24352 22704 24404
rect 7656 24284 7708 24336
rect 8944 24284 8996 24336
rect 14372 24284 14424 24336
rect 17500 24327 17552 24336
rect 7104 24216 7156 24268
rect 5264 24148 5316 24200
rect 5172 24080 5224 24132
rect 7656 24148 7708 24200
rect 7840 24080 7892 24132
rect 9496 24216 9548 24268
rect 9956 24216 10008 24268
rect 13176 24216 13228 24268
rect 15476 24216 15528 24268
rect 17500 24293 17509 24327
rect 17509 24293 17543 24327
rect 17543 24293 17552 24327
rect 17500 24284 17552 24293
rect 16120 24216 16172 24268
rect 19524 24216 19576 24268
rect 15200 24148 15252 24200
rect 15292 24148 15344 24200
rect 12808 24080 12860 24132
rect 12992 24080 13044 24132
rect 13912 24080 13964 24132
rect 17408 24080 17460 24132
rect 17684 24123 17736 24132
rect 17684 24089 17693 24123
rect 17693 24089 17727 24123
rect 17727 24089 17736 24123
rect 17684 24080 17736 24089
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 9680 24012 9732 24064
rect 14004 24012 14056 24064
rect 16212 24012 16264 24064
rect 22100 24259 22152 24268
rect 22100 24225 22109 24259
rect 22109 24225 22143 24259
rect 22143 24225 22152 24259
rect 22100 24216 22152 24225
rect 22468 24216 22520 24268
rect 22928 24259 22980 24268
rect 22928 24225 22937 24259
rect 22937 24225 22971 24259
rect 22971 24225 22980 24259
rect 22928 24216 22980 24225
rect 26424 24352 26476 24404
rect 26700 24284 26752 24336
rect 26056 24191 26108 24200
rect 26056 24157 26065 24191
rect 26065 24157 26099 24191
rect 26099 24157 26108 24191
rect 26056 24148 26108 24157
rect 22100 24080 22152 24132
rect 22192 24012 22244 24064
rect 23020 24012 23072 24064
rect 5536 23910 5588 23962
rect 5600 23910 5652 23962
rect 5664 23910 5716 23962
rect 5728 23910 5780 23962
rect 14644 23910 14696 23962
rect 14708 23910 14760 23962
rect 14772 23910 14824 23962
rect 14836 23910 14888 23962
rect 23752 23910 23804 23962
rect 23816 23910 23868 23962
rect 23880 23910 23932 23962
rect 23944 23910 23996 23962
rect 2872 23808 2924 23860
rect 6920 23808 6972 23860
rect 7564 23808 7616 23860
rect 9956 23783 10008 23792
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 9956 23749 9965 23783
rect 9965 23749 9999 23783
rect 9999 23749 10008 23783
rect 9956 23740 10008 23749
rect 16212 23740 16264 23792
rect 1584 23604 1636 23656
rect 4528 23604 4580 23656
rect 7472 23604 7524 23656
rect 7564 23647 7616 23656
rect 7564 23613 7573 23647
rect 7573 23613 7607 23647
rect 7607 23613 7616 23647
rect 9404 23647 9456 23656
rect 7564 23604 7616 23613
rect 9404 23613 9413 23647
rect 9413 23613 9447 23647
rect 9447 23613 9456 23647
rect 9404 23604 9456 23613
rect 9680 23647 9732 23656
rect 3056 23536 3108 23588
rect 9680 23613 9689 23647
rect 9689 23613 9723 23647
rect 9723 23613 9732 23647
rect 9680 23604 9732 23613
rect 10508 23672 10560 23724
rect 10784 23715 10836 23724
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 11336 23672 11388 23724
rect 13360 23672 13412 23724
rect 10416 23647 10468 23656
rect 10416 23613 10425 23647
rect 10425 23613 10459 23647
rect 10459 23613 10468 23647
rect 10416 23604 10468 23613
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 10968 23647 11020 23656
rect 10968 23613 10977 23647
rect 10977 23613 11011 23647
rect 11011 23613 11020 23647
rect 10968 23604 11020 23613
rect 13728 23672 13780 23724
rect 15476 23672 15528 23724
rect 14096 23647 14148 23656
rect 14096 23613 14105 23647
rect 14105 23613 14139 23647
rect 14139 23613 14148 23647
rect 14096 23604 14148 23613
rect 15200 23604 15252 23656
rect 17684 23808 17736 23860
rect 19524 23851 19576 23860
rect 19524 23817 19533 23851
rect 19533 23817 19567 23851
rect 19567 23817 19576 23851
rect 19524 23808 19576 23817
rect 23204 23740 23256 23792
rect 22652 23672 22704 23724
rect 22744 23647 22796 23656
rect 3884 23511 3936 23520
rect 3884 23477 3893 23511
rect 3893 23477 3927 23511
rect 3927 23477 3936 23511
rect 3884 23468 3936 23477
rect 6736 23468 6788 23520
rect 10784 23536 10836 23588
rect 13176 23536 13228 23588
rect 15292 23579 15344 23588
rect 15292 23545 15301 23579
rect 15301 23545 15335 23579
rect 15335 23545 15344 23579
rect 15292 23536 15344 23545
rect 17224 23536 17276 23588
rect 22744 23613 22753 23647
rect 22753 23613 22787 23647
rect 22787 23613 22796 23647
rect 22744 23604 22796 23613
rect 23940 23647 23992 23656
rect 18420 23579 18472 23588
rect 18420 23545 18454 23579
rect 18454 23545 18472 23579
rect 18420 23536 18472 23545
rect 20628 23536 20680 23588
rect 21548 23536 21600 23588
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 26424 23672 26476 23724
rect 26148 23647 26200 23656
rect 26148 23613 26157 23647
rect 26157 23613 26191 23647
rect 26191 23613 26200 23647
rect 26148 23604 26200 23613
rect 26608 23604 26660 23656
rect 24216 23579 24268 23588
rect 24216 23545 24250 23579
rect 24250 23545 24268 23579
rect 24216 23536 24268 23545
rect 12992 23468 13044 23520
rect 13636 23511 13688 23520
rect 13636 23477 13645 23511
rect 13645 23477 13679 23511
rect 13679 23477 13688 23511
rect 13636 23468 13688 23477
rect 14188 23511 14240 23520
rect 14188 23477 14197 23511
rect 14197 23477 14231 23511
rect 14231 23477 14240 23511
rect 14188 23468 14240 23477
rect 15016 23468 15068 23520
rect 15844 23468 15896 23520
rect 17960 23468 18012 23520
rect 21272 23468 21324 23520
rect 21456 23511 21508 23520
rect 21456 23477 21465 23511
rect 21465 23477 21499 23511
rect 21499 23477 21508 23511
rect 21456 23468 21508 23477
rect 23572 23468 23624 23520
rect 25320 23511 25372 23520
rect 25320 23477 25329 23511
rect 25329 23477 25363 23511
rect 25363 23477 25372 23511
rect 25320 23468 25372 23477
rect 26148 23468 26200 23520
rect 26700 23511 26752 23520
rect 26700 23477 26709 23511
rect 26709 23477 26743 23511
rect 26743 23477 26752 23511
rect 26700 23468 26752 23477
rect 10090 23366 10142 23418
rect 10154 23366 10206 23418
rect 10218 23366 10270 23418
rect 10282 23366 10334 23418
rect 19198 23366 19250 23418
rect 19262 23366 19314 23418
rect 19326 23366 19378 23418
rect 19390 23366 19442 23418
rect 3056 23307 3108 23316
rect 3056 23273 3065 23307
rect 3065 23273 3099 23307
rect 3099 23273 3108 23307
rect 3056 23264 3108 23273
rect 5264 23264 5316 23316
rect 1860 23239 1912 23248
rect 1860 23205 1869 23239
rect 1869 23205 1903 23239
rect 1903 23205 1912 23239
rect 1860 23196 1912 23205
rect 3884 23196 3936 23248
rect 10416 23264 10468 23316
rect 10968 23264 11020 23316
rect 15108 23264 15160 23316
rect 17316 23264 17368 23316
rect 18420 23307 18472 23316
rect 18420 23273 18429 23307
rect 18429 23273 18463 23307
rect 18463 23273 18472 23307
rect 18420 23264 18472 23273
rect 18696 23264 18748 23316
rect 21180 23264 21232 23316
rect 22744 23264 22796 23316
rect 26148 23264 26200 23316
rect 2504 23171 2556 23180
rect 2504 23137 2513 23171
rect 2513 23137 2547 23171
rect 2547 23137 2556 23171
rect 2504 23128 2556 23137
rect 2596 23128 2648 23180
rect 3148 23128 3200 23180
rect 6644 23171 6696 23180
rect 6644 23137 6653 23171
rect 6653 23137 6687 23171
rect 6687 23137 6696 23171
rect 6644 23128 6696 23137
rect 14464 23196 14516 23248
rect 6000 22992 6052 23044
rect 9680 23128 9732 23180
rect 11980 23128 12032 23180
rect 12992 23171 13044 23180
rect 12992 23137 13001 23171
rect 13001 23137 13035 23171
rect 13035 23137 13044 23171
rect 12992 23128 13044 23137
rect 13084 23128 13136 23180
rect 13452 23171 13504 23180
rect 13452 23137 13461 23171
rect 13461 23137 13495 23171
rect 13495 23137 13504 23171
rect 13452 23128 13504 23137
rect 14188 23128 14240 23180
rect 14832 23171 14884 23180
rect 14832 23137 14841 23171
rect 14841 23137 14875 23171
rect 14875 23137 14884 23171
rect 14832 23128 14884 23137
rect 15660 23128 15712 23180
rect 16212 23171 16264 23180
rect 16212 23137 16221 23171
rect 16221 23137 16255 23171
rect 16255 23137 16264 23171
rect 16212 23128 16264 23137
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 17868 23171 17920 23180
rect 10968 23060 11020 23112
rect 15016 23060 15068 23112
rect 11060 22992 11112 23044
rect 13544 23035 13596 23044
rect 13544 23001 13553 23035
rect 13553 23001 13587 23035
rect 13587 23001 13596 23035
rect 13544 22992 13596 23001
rect 16028 22992 16080 23044
rect 17224 23035 17276 23044
rect 17224 23001 17233 23035
rect 17233 23001 17267 23035
rect 17267 23001 17276 23035
rect 17224 22992 17276 23001
rect 1952 22967 2004 22976
rect 1952 22933 1961 22967
rect 1961 22933 1995 22967
rect 1995 22933 2004 22967
rect 1952 22924 2004 22933
rect 6920 22924 6972 22976
rect 8208 22924 8260 22976
rect 10508 22924 10560 22976
rect 10876 22924 10928 22976
rect 12072 22924 12124 22976
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 18788 23196 18840 23248
rect 24308 23196 24360 23248
rect 26700 23196 26752 23248
rect 18236 23171 18288 23180
rect 18236 23137 18245 23171
rect 18245 23137 18279 23171
rect 18279 23137 18288 23171
rect 18236 23128 18288 23137
rect 18880 23128 18932 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 18696 23060 18748 23112
rect 20444 23171 20496 23180
rect 20444 23137 20453 23171
rect 20453 23137 20487 23171
rect 20487 23137 20496 23171
rect 20444 23128 20496 23137
rect 21640 23128 21692 23180
rect 21456 23060 21508 23112
rect 21548 23103 21600 23112
rect 21548 23069 21557 23103
rect 21557 23069 21591 23103
rect 21591 23069 21600 23103
rect 21548 23060 21600 23069
rect 18144 22992 18196 23044
rect 19524 22992 19576 23044
rect 20628 23035 20680 23044
rect 20628 23001 20637 23035
rect 20637 23001 20671 23035
rect 20671 23001 20680 23035
rect 20628 22992 20680 23001
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 21364 22924 21416 22976
rect 24124 23128 24176 23180
rect 26056 23103 26108 23112
rect 23480 22992 23532 23044
rect 23940 22992 23992 23044
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 24308 22924 24360 22976
rect 25320 22924 25372 22976
rect 5536 22822 5588 22874
rect 5600 22822 5652 22874
rect 5664 22822 5716 22874
rect 5728 22822 5780 22874
rect 14644 22822 14696 22874
rect 14708 22822 14760 22874
rect 14772 22822 14824 22874
rect 14836 22822 14888 22874
rect 23752 22822 23804 22874
rect 23816 22822 23868 22874
rect 23880 22822 23932 22874
rect 23944 22822 23996 22874
rect 5172 22720 5224 22772
rect 10416 22763 10468 22772
rect 10416 22729 10425 22763
rect 10425 22729 10459 22763
rect 10459 22729 10468 22763
rect 10416 22720 10468 22729
rect 10600 22720 10652 22772
rect 14096 22720 14148 22772
rect 1952 22652 2004 22704
rect 5264 22516 5316 22568
rect 6276 22516 6328 22568
rect 6828 22559 6880 22568
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 7380 22584 7432 22636
rect 9680 22584 9732 22636
rect 11060 22652 11112 22704
rect 2044 22491 2096 22500
rect 2044 22457 2053 22491
rect 2053 22457 2087 22491
rect 2087 22457 2096 22491
rect 2044 22448 2096 22457
rect 7288 22516 7340 22568
rect 7564 22516 7616 22568
rect 8944 22559 8996 22568
rect 8944 22525 8953 22559
rect 8953 22525 8987 22559
rect 8987 22525 8996 22559
rect 8944 22516 8996 22525
rect 9128 22516 9180 22568
rect 10232 22559 10284 22568
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 12256 22584 12308 22636
rect 13820 22652 13872 22704
rect 15016 22720 15068 22772
rect 7104 22491 7156 22500
rect 7104 22457 7113 22491
rect 7113 22457 7147 22491
rect 7147 22457 7156 22491
rect 7104 22448 7156 22457
rect 7012 22380 7064 22432
rect 9588 22448 9640 22500
rect 7380 22423 7432 22432
rect 7380 22389 7389 22423
rect 7389 22389 7423 22423
rect 7423 22389 7432 22423
rect 7380 22380 7432 22389
rect 8852 22380 8904 22432
rect 9220 22380 9272 22432
rect 10600 22448 10652 22500
rect 11612 22516 11664 22568
rect 12072 22559 12124 22568
rect 12072 22525 12081 22559
rect 12081 22525 12115 22559
rect 12115 22525 12124 22559
rect 12072 22516 12124 22525
rect 12716 22516 12768 22568
rect 11152 22380 11204 22432
rect 13636 22448 13688 22500
rect 15476 22652 15528 22704
rect 16396 22695 16448 22704
rect 16396 22661 16405 22695
rect 16405 22661 16439 22695
rect 16439 22661 16448 22695
rect 16396 22652 16448 22661
rect 15476 22559 15528 22568
rect 15476 22525 15485 22559
rect 15485 22525 15519 22559
rect 15519 22525 15528 22559
rect 17868 22584 17920 22636
rect 17316 22559 17368 22568
rect 15476 22516 15528 22525
rect 17316 22525 17325 22559
rect 17325 22525 17359 22559
rect 17359 22525 17368 22559
rect 17316 22516 17368 22525
rect 17592 22559 17644 22568
rect 17592 22525 17601 22559
rect 17601 22525 17635 22559
rect 17635 22525 17644 22559
rect 17592 22516 17644 22525
rect 17684 22559 17736 22568
rect 17684 22525 17693 22559
rect 17693 22525 17727 22559
rect 17727 22525 17736 22559
rect 17684 22516 17736 22525
rect 18236 22516 18288 22568
rect 18328 22516 18380 22568
rect 20536 22584 20588 22636
rect 22192 22652 22244 22704
rect 23296 22652 23348 22704
rect 23940 22652 23992 22704
rect 21916 22584 21968 22636
rect 20076 22516 20128 22568
rect 21364 22559 21416 22568
rect 16120 22448 16172 22500
rect 17408 22448 17460 22500
rect 18420 22448 18472 22500
rect 19156 22448 19208 22500
rect 19984 22448 20036 22500
rect 17868 22423 17920 22432
rect 17868 22389 17877 22423
rect 17877 22389 17911 22423
rect 17911 22389 17920 22423
rect 17868 22380 17920 22389
rect 18052 22380 18104 22432
rect 18788 22380 18840 22432
rect 19800 22380 19852 22432
rect 20628 22380 20680 22432
rect 21364 22525 21373 22559
rect 21373 22525 21407 22559
rect 21407 22525 21416 22559
rect 21364 22516 21416 22525
rect 21456 22559 21508 22568
rect 21456 22525 21489 22559
rect 21489 22525 21508 22559
rect 21456 22516 21508 22525
rect 21640 22516 21692 22568
rect 23480 22584 23532 22636
rect 21272 22491 21324 22500
rect 21272 22457 21281 22491
rect 21281 22457 21315 22491
rect 21315 22457 21324 22491
rect 21272 22448 21324 22457
rect 24584 22516 24636 22568
rect 26148 22516 26200 22568
rect 26792 22516 26844 22568
rect 22652 22448 22704 22500
rect 22560 22380 22612 22432
rect 25780 22448 25832 22500
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 25412 22423 25464 22432
rect 25412 22389 25421 22423
rect 25421 22389 25455 22423
rect 25455 22389 25464 22423
rect 25412 22380 25464 22389
rect 10090 22278 10142 22330
rect 10154 22278 10206 22330
rect 10218 22278 10270 22330
rect 10282 22278 10334 22330
rect 19198 22278 19250 22330
rect 19262 22278 19314 22330
rect 19326 22278 19378 22330
rect 19390 22278 19442 22330
rect 5172 22040 5224 22092
rect 6644 22176 6696 22228
rect 6828 22176 6880 22228
rect 6920 22176 6972 22228
rect 7288 22176 7340 22228
rect 11980 22219 12032 22228
rect 11980 22185 11989 22219
rect 11989 22185 12023 22219
rect 12023 22185 12032 22219
rect 11980 22176 12032 22185
rect 12716 22176 12768 22228
rect 13452 22176 13504 22228
rect 17040 22176 17092 22228
rect 17592 22219 17644 22228
rect 17592 22185 17601 22219
rect 17601 22185 17635 22219
rect 17635 22185 17644 22219
rect 17592 22176 17644 22185
rect 18420 22176 18472 22228
rect 22652 22176 22704 22228
rect 22928 22176 22980 22228
rect 6460 22108 6512 22160
rect 7564 22040 7616 22092
rect 6736 21972 6788 22024
rect 7196 21972 7248 22024
rect 9128 22040 9180 22092
rect 9588 22040 9640 22092
rect 10692 22108 10744 22160
rect 12072 22108 12124 22160
rect 10048 22040 10100 22092
rect 10600 22040 10652 22092
rect 10876 22040 10928 22092
rect 11428 22083 11480 22092
rect 11428 22049 11437 22083
rect 11437 22049 11471 22083
rect 11471 22049 11480 22083
rect 11428 22040 11480 22049
rect 15936 22108 15988 22160
rect 9680 21904 9732 21956
rect 9772 21904 9824 21956
rect 10692 21904 10744 21956
rect 11704 21972 11756 22024
rect 12992 22040 13044 22092
rect 15292 22040 15344 22092
rect 15844 22040 15896 22092
rect 17868 22040 17920 22092
rect 19248 22108 19300 22160
rect 20536 22108 20588 22160
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 17408 21972 17460 22024
rect 19800 21972 19852 22024
rect 13268 21904 13320 21956
rect 18328 21904 18380 21956
rect 18972 21904 19024 21956
rect 19248 21904 19300 21956
rect 20260 22083 20312 22092
rect 20260 22049 20269 22083
rect 20269 22049 20303 22083
rect 20303 22049 20312 22083
rect 20260 22040 20312 22049
rect 20444 22040 20496 22092
rect 21456 22108 21508 22160
rect 21916 22108 21968 22160
rect 23112 22108 23164 22160
rect 24400 22176 24452 22228
rect 25412 22176 25464 22228
rect 25780 22219 25832 22228
rect 25780 22185 25789 22219
rect 25789 22185 25823 22219
rect 25823 22185 25832 22219
rect 25780 22176 25832 22185
rect 21548 22040 21600 22092
rect 23480 22040 23532 22092
rect 23572 22040 23624 22092
rect 23848 22083 23900 22092
rect 23848 22049 23857 22083
rect 23857 22049 23891 22083
rect 23891 22049 23900 22083
rect 23848 22040 23900 22049
rect 23940 22083 23992 22092
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 24768 22040 24820 22092
rect 25228 22083 25280 22092
rect 25228 22049 25237 22083
rect 25237 22049 25271 22083
rect 25271 22049 25280 22083
rect 25228 22040 25280 22049
rect 27252 22108 27304 22160
rect 27528 22151 27580 22160
rect 27528 22117 27537 22151
rect 27537 22117 27571 22151
rect 27571 22117 27580 22151
rect 27528 22108 27580 22117
rect 25688 22040 25740 22092
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 20076 21904 20128 21956
rect 20168 21904 20220 21956
rect 23388 21904 23440 21956
rect 6552 21836 6604 21888
rect 6736 21836 6788 21888
rect 7196 21836 7248 21888
rect 8116 21836 8168 21888
rect 9956 21836 10008 21888
rect 10508 21836 10560 21888
rect 11152 21836 11204 21888
rect 11704 21836 11756 21888
rect 12808 21836 12860 21888
rect 12992 21836 13044 21888
rect 13452 21836 13504 21888
rect 13728 21836 13780 21888
rect 15200 21836 15252 21888
rect 15292 21836 15344 21888
rect 15476 21836 15528 21888
rect 17316 21836 17368 21888
rect 18696 21836 18748 21888
rect 20536 21879 20588 21888
rect 20536 21845 20545 21879
rect 20545 21845 20579 21879
rect 20579 21845 20588 21879
rect 20536 21836 20588 21845
rect 22560 21836 22612 21888
rect 23572 21836 23624 21888
rect 23848 21904 23900 21956
rect 25412 21904 25464 21956
rect 27620 21879 27672 21888
rect 27620 21845 27629 21879
rect 27629 21845 27663 21879
rect 27663 21845 27672 21879
rect 27620 21836 27672 21845
rect 5536 21734 5588 21786
rect 5600 21734 5652 21786
rect 5664 21734 5716 21786
rect 5728 21734 5780 21786
rect 14644 21734 14696 21786
rect 14708 21734 14760 21786
rect 14772 21734 14824 21786
rect 14836 21734 14888 21786
rect 23752 21734 23804 21786
rect 23816 21734 23868 21786
rect 23880 21734 23932 21786
rect 23944 21734 23996 21786
rect 6736 21632 6788 21684
rect 7104 21632 7156 21684
rect 8208 21675 8260 21684
rect 8208 21641 8217 21675
rect 8217 21641 8251 21675
rect 8251 21641 8260 21675
rect 8208 21632 8260 21641
rect 8484 21632 8536 21684
rect 3884 21564 3936 21616
rect 4712 21564 4764 21616
rect 5724 21564 5776 21616
rect 8944 21564 8996 21616
rect 9680 21564 9732 21616
rect 10692 21632 10744 21684
rect 12348 21632 12400 21684
rect 14832 21564 14884 21616
rect 16120 21564 16172 21616
rect 16396 21564 16448 21616
rect 1676 21471 1728 21480
rect 1676 21437 1685 21471
rect 1685 21437 1719 21471
rect 1719 21437 1728 21471
rect 1676 21428 1728 21437
rect 2136 21471 2188 21480
rect 2136 21437 2145 21471
rect 2145 21437 2179 21471
rect 2179 21437 2188 21471
rect 2136 21428 2188 21437
rect 3608 21428 3660 21480
rect 3332 21360 3384 21412
rect 5448 21428 5500 21480
rect 12900 21496 12952 21548
rect 13636 21496 13688 21548
rect 15016 21496 15068 21548
rect 18236 21632 18288 21684
rect 18420 21632 18472 21684
rect 19248 21632 19300 21684
rect 23020 21675 23072 21684
rect 17040 21564 17092 21616
rect 17500 21564 17552 21616
rect 17592 21564 17644 21616
rect 5724 21471 5776 21480
rect 5724 21437 5733 21471
rect 5733 21437 5767 21471
rect 5767 21437 5776 21471
rect 5724 21428 5776 21437
rect 5816 21428 5868 21480
rect 6368 21428 6420 21480
rect 6644 21428 6696 21480
rect 6920 21428 6972 21480
rect 7380 21428 7432 21480
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 9220 21471 9272 21480
rect 7564 21360 7616 21412
rect 8300 21360 8352 21412
rect 9220 21437 9229 21471
rect 9229 21437 9263 21471
rect 9263 21437 9272 21471
rect 9220 21428 9272 21437
rect 9680 21471 9732 21480
rect 9680 21437 9689 21471
rect 9689 21437 9723 21471
rect 9723 21437 9732 21471
rect 9680 21428 9732 21437
rect 9956 21471 10008 21480
rect 9956 21437 9990 21471
rect 9990 21437 10008 21471
rect 9956 21428 10008 21437
rect 12348 21428 12400 21480
rect 12716 21428 12768 21480
rect 13728 21428 13780 21480
rect 14188 21428 14240 21480
rect 15292 21428 15344 21480
rect 15476 21428 15528 21480
rect 17040 21428 17092 21480
rect 3792 21292 3844 21344
rect 4160 21335 4212 21344
rect 4160 21301 4169 21335
rect 4169 21301 4203 21335
rect 4203 21301 4212 21335
rect 4160 21292 4212 21301
rect 4896 21292 4948 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 9312 21292 9364 21344
rect 9404 21292 9456 21344
rect 10784 21292 10836 21344
rect 12624 21292 12676 21344
rect 13268 21292 13320 21344
rect 13728 21292 13780 21344
rect 15936 21360 15988 21412
rect 18236 21428 18288 21480
rect 18604 21428 18656 21480
rect 18972 21564 19024 21616
rect 20904 21496 20956 21548
rect 18972 21428 19024 21480
rect 19156 21428 19208 21480
rect 20536 21428 20588 21480
rect 20628 21428 20680 21480
rect 22652 21428 22704 21480
rect 23020 21641 23029 21675
rect 23029 21641 23063 21675
rect 23063 21641 23072 21675
rect 23020 21632 23072 21641
rect 24216 21675 24268 21684
rect 24216 21641 24225 21675
rect 24225 21641 24259 21675
rect 24259 21641 24268 21675
rect 24216 21632 24268 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 25412 21675 25464 21684
rect 25412 21641 25421 21675
rect 25421 21641 25455 21675
rect 25455 21641 25464 21675
rect 25412 21632 25464 21641
rect 23204 21564 23256 21616
rect 23664 21564 23716 21616
rect 23940 21564 23992 21616
rect 25688 21564 25740 21616
rect 24584 21496 24636 21548
rect 23572 21428 23624 21480
rect 23940 21471 23992 21480
rect 23940 21437 23949 21471
rect 23949 21437 23983 21471
rect 23983 21437 23992 21471
rect 23940 21428 23992 21437
rect 24308 21428 24360 21480
rect 24492 21428 24544 21480
rect 25596 21428 25648 21480
rect 14280 21292 14332 21344
rect 15108 21292 15160 21344
rect 15200 21292 15252 21344
rect 16120 21292 16172 21344
rect 18052 21292 18104 21344
rect 18604 21292 18656 21344
rect 19524 21292 19576 21344
rect 20260 21292 20312 21344
rect 23112 21292 23164 21344
rect 24216 21360 24268 21412
rect 24768 21360 24820 21412
rect 25228 21360 25280 21412
rect 25688 21292 25740 21344
rect 25780 21292 25832 21344
rect 26976 21360 27028 21412
rect 26516 21335 26568 21344
rect 26516 21301 26525 21335
rect 26525 21301 26559 21335
rect 26559 21301 26568 21335
rect 26516 21292 26568 21301
rect 10090 21190 10142 21242
rect 10154 21190 10206 21242
rect 10218 21190 10270 21242
rect 10282 21190 10334 21242
rect 19198 21190 19250 21242
rect 19262 21190 19314 21242
rect 19326 21190 19378 21242
rect 19390 21190 19442 21242
rect 1952 21131 2004 21140
rect 1952 21097 1961 21131
rect 1961 21097 1995 21131
rect 1995 21097 2004 21131
rect 1952 21088 2004 21097
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 4160 21020 4212 21072
rect 1860 20995 1912 21004
rect 1860 20961 1869 20995
rect 1869 20961 1903 20995
rect 1903 20961 1912 20995
rect 1860 20952 1912 20961
rect 3884 20952 3936 21004
rect 6000 21088 6052 21140
rect 6368 21088 6420 21140
rect 9404 21088 9456 21140
rect 9680 21088 9732 21140
rect 10784 21088 10836 21140
rect 10876 21088 10928 21140
rect 4896 20995 4948 21004
rect 4896 20961 4905 20995
rect 4905 20961 4939 20995
rect 4939 20961 4948 20995
rect 4896 20952 4948 20961
rect 5816 21020 5868 21072
rect 5908 21020 5960 21072
rect 6736 21020 6788 21072
rect 5264 20995 5316 21004
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 7932 20952 7984 21004
rect 3056 20884 3108 20936
rect 5816 20884 5868 20936
rect 4252 20748 4304 20800
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 8300 20952 8352 20961
rect 8668 20952 8720 21004
rect 9496 20995 9548 21004
rect 9496 20961 9505 20995
rect 9505 20961 9539 20995
rect 9539 20961 9548 20995
rect 9496 20952 9548 20961
rect 10416 21020 10468 21072
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 13360 20952 13412 21004
rect 15936 21020 15988 21072
rect 17132 21020 17184 21072
rect 17684 21020 17736 21072
rect 20076 21088 20128 21140
rect 22468 21088 22520 21140
rect 22652 21131 22704 21140
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 20996 21020 21048 21072
rect 23020 21020 23072 21072
rect 14464 20952 14516 21004
rect 14832 20952 14884 21004
rect 15200 20952 15252 21004
rect 15476 20952 15528 21004
rect 17040 20952 17092 21004
rect 8300 20816 8352 20868
rect 13636 20884 13688 20936
rect 13728 20884 13780 20936
rect 15108 20927 15160 20936
rect 14832 20816 14884 20868
rect 15108 20893 15117 20927
rect 15117 20893 15151 20927
rect 15151 20893 15160 20927
rect 15108 20884 15160 20893
rect 17316 20884 17368 20936
rect 18236 20995 18288 21004
rect 18236 20961 18245 20995
rect 18245 20961 18279 20995
rect 18279 20961 18288 20995
rect 18512 20995 18564 21004
rect 18236 20952 18288 20961
rect 18512 20961 18521 20995
rect 18521 20961 18555 20995
rect 18555 20961 18564 20995
rect 18512 20952 18564 20961
rect 18696 20952 18748 21004
rect 19616 20884 19668 20936
rect 19984 20952 20036 21004
rect 20444 20952 20496 21004
rect 20720 20995 20772 21004
rect 20720 20961 20729 20995
rect 20729 20961 20763 20995
rect 20763 20961 20772 20995
rect 20720 20952 20772 20961
rect 21824 20995 21876 21004
rect 21824 20961 21833 20995
rect 21833 20961 21867 20995
rect 21867 20961 21876 20995
rect 21824 20952 21876 20961
rect 22560 20995 22612 21004
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 24400 21088 24452 21140
rect 24584 20952 24636 21004
rect 25228 20952 25280 21004
rect 15568 20816 15620 20868
rect 18420 20859 18472 20868
rect 6184 20748 6236 20800
rect 7564 20748 7616 20800
rect 8392 20748 8444 20800
rect 8944 20748 8996 20800
rect 10692 20748 10744 20800
rect 12256 20748 12308 20800
rect 14188 20748 14240 20800
rect 15384 20791 15436 20800
rect 15384 20757 15393 20791
rect 15393 20757 15427 20791
rect 15427 20757 15436 20791
rect 15384 20748 15436 20757
rect 15844 20748 15896 20800
rect 17776 20748 17828 20800
rect 18420 20825 18429 20859
rect 18429 20825 18463 20859
rect 18463 20825 18472 20859
rect 18420 20816 18472 20825
rect 19340 20816 19392 20868
rect 21272 20816 21324 20868
rect 22468 20816 22520 20868
rect 25596 20995 25648 21004
rect 25596 20961 25605 20995
rect 25605 20961 25639 20995
rect 25639 20961 25648 20995
rect 25596 20952 25648 20961
rect 25688 20995 25740 21004
rect 25688 20961 25697 20995
rect 25697 20961 25731 20995
rect 25731 20961 25740 20995
rect 25688 20952 25740 20961
rect 26056 20952 26108 21004
rect 27068 20952 27120 21004
rect 27344 20952 27396 21004
rect 23480 20748 23532 20800
rect 24124 20748 24176 20800
rect 27344 20748 27396 20800
rect 5536 20646 5588 20698
rect 5600 20646 5652 20698
rect 5664 20646 5716 20698
rect 5728 20646 5780 20698
rect 14644 20646 14696 20698
rect 14708 20646 14760 20698
rect 14772 20646 14824 20698
rect 14836 20646 14888 20698
rect 23752 20646 23804 20698
rect 23816 20646 23868 20698
rect 23880 20646 23932 20698
rect 23944 20646 23996 20698
rect 5264 20544 5316 20596
rect 5908 20544 5960 20596
rect 7104 20544 7156 20596
rect 8576 20587 8628 20596
rect 8576 20553 8585 20587
rect 8585 20553 8619 20587
rect 8619 20553 8628 20587
rect 8576 20544 8628 20553
rect 9496 20544 9548 20596
rect 12348 20544 12400 20596
rect 14188 20544 14240 20596
rect 15108 20544 15160 20596
rect 18420 20544 18472 20596
rect 19616 20587 19668 20596
rect 19616 20553 19625 20587
rect 19625 20553 19659 20587
rect 19659 20553 19668 20587
rect 19616 20544 19668 20553
rect 10968 20476 11020 20528
rect 13268 20476 13320 20528
rect 6644 20408 6696 20460
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 2872 20272 2924 20324
rect 2688 20204 2740 20256
rect 3608 20340 3660 20392
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 10508 20408 10560 20460
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 25504 20544 25556 20596
rect 24768 20476 24820 20528
rect 15752 20451 15804 20460
rect 14096 20408 14148 20417
rect 10416 20340 10468 20392
rect 5816 20272 5868 20324
rect 7472 20315 7524 20324
rect 7472 20281 7506 20315
rect 7506 20281 7524 20315
rect 7472 20272 7524 20281
rect 10508 20272 10560 20324
rect 11060 20340 11112 20392
rect 11244 20340 11296 20392
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 13728 20315 13780 20324
rect 5540 20204 5592 20256
rect 13728 20281 13737 20315
rect 13737 20281 13771 20315
rect 13771 20281 13780 20315
rect 13728 20272 13780 20281
rect 15108 20340 15160 20392
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 15936 20340 15988 20392
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 18236 20340 18288 20392
rect 18696 20340 18748 20392
rect 18972 20408 19024 20460
rect 23480 20451 23532 20460
rect 19340 20340 19392 20392
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 17224 20272 17276 20324
rect 20076 20272 20128 20324
rect 20352 20272 20404 20324
rect 14280 20204 14332 20256
rect 18788 20204 18840 20256
rect 21824 20272 21876 20324
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 23480 20408 23532 20417
rect 23112 20383 23164 20392
rect 23112 20349 23121 20383
rect 23121 20349 23155 20383
rect 23155 20349 23164 20383
rect 23112 20340 23164 20349
rect 23296 20340 23348 20392
rect 24124 20383 24176 20392
rect 23388 20272 23440 20324
rect 24124 20349 24133 20383
rect 24133 20349 24167 20383
rect 24167 20349 24176 20383
rect 24124 20340 24176 20349
rect 24860 20383 24912 20392
rect 24860 20349 24869 20383
rect 24869 20349 24903 20383
rect 24903 20349 24912 20383
rect 24860 20340 24912 20349
rect 25136 20272 25188 20324
rect 26516 20340 26568 20392
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 25780 20204 25832 20256
rect 26976 20204 27028 20256
rect 10090 20102 10142 20154
rect 10154 20102 10206 20154
rect 10218 20102 10270 20154
rect 10282 20102 10334 20154
rect 19198 20102 19250 20154
rect 19262 20102 19314 20154
rect 19326 20102 19378 20154
rect 19390 20102 19442 20154
rect 2872 20000 2924 20052
rect 5816 20043 5868 20052
rect 5816 20009 5825 20043
rect 5825 20009 5859 20043
rect 5859 20009 5868 20043
rect 5816 20000 5868 20009
rect 6276 20043 6328 20052
rect 6276 20009 6285 20043
rect 6285 20009 6319 20043
rect 6319 20009 6328 20043
rect 6276 20000 6328 20009
rect 6736 20000 6788 20052
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 9680 20000 9732 20052
rect 10508 20000 10560 20052
rect 3056 19932 3108 19984
rect 5540 19975 5592 19984
rect 2228 19864 2280 19916
rect 2412 19907 2464 19916
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2412 19864 2464 19873
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 3976 19864 4028 19916
rect 5540 19941 5549 19975
rect 5549 19941 5583 19975
rect 5583 19941 5592 19975
rect 5540 19932 5592 19941
rect 5908 19932 5960 19984
rect 5448 19907 5500 19916
rect 1676 19796 1728 19848
rect 5448 19873 5457 19907
rect 5457 19873 5491 19907
rect 5491 19873 5500 19907
rect 5448 19864 5500 19873
rect 6000 19864 6052 19916
rect 6552 19932 6604 19984
rect 7012 19932 7064 19984
rect 8576 19932 8628 19984
rect 6920 19907 6972 19916
rect 6368 19796 6420 19848
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 7472 19864 7524 19916
rect 8208 19907 8260 19916
rect 8208 19873 8217 19907
rect 8217 19873 8251 19907
rect 8251 19873 8260 19907
rect 8208 19864 8260 19873
rect 8392 19864 8444 19916
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 10416 19907 10468 19916
rect 10416 19873 10425 19907
rect 10425 19873 10459 19907
rect 10459 19873 10468 19907
rect 10416 19864 10468 19873
rect 10692 19907 10744 19916
rect 10692 19873 10701 19907
rect 10701 19873 10735 19907
rect 10735 19873 10744 19907
rect 10692 19864 10744 19873
rect 11336 20000 11388 20052
rect 13084 20000 13136 20052
rect 15384 20000 15436 20052
rect 1952 19771 2004 19780
rect 1952 19737 1961 19771
rect 1961 19737 1995 19771
rect 1995 19737 2004 19771
rect 1952 19728 2004 19737
rect 7840 19796 7892 19848
rect 13360 19932 13412 19984
rect 11888 19907 11940 19916
rect 11888 19873 11897 19907
rect 11897 19873 11931 19907
rect 11931 19873 11940 19907
rect 11888 19864 11940 19873
rect 13728 19864 13780 19916
rect 18328 19932 18380 19984
rect 18696 19932 18748 19984
rect 21824 20000 21876 20052
rect 22652 20000 22704 20052
rect 27068 20000 27120 20052
rect 21180 19932 21232 19984
rect 22928 19932 22980 19984
rect 23572 19932 23624 19984
rect 24124 19975 24176 19984
rect 24124 19941 24133 19975
rect 24133 19941 24167 19975
rect 24167 19941 24176 19975
rect 24124 19932 24176 19941
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 15292 19864 15344 19916
rect 16212 19907 16264 19916
rect 16212 19873 16221 19907
rect 16221 19873 16255 19907
rect 16255 19873 16264 19907
rect 16212 19864 16264 19873
rect 17316 19864 17368 19916
rect 18420 19864 18472 19916
rect 18972 19864 19024 19916
rect 22744 19864 22796 19916
rect 15476 19839 15528 19848
rect 13452 19796 13504 19805
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 19800 19796 19852 19848
rect 23204 19907 23256 19916
rect 23204 19873 23213 19907
rect 23213 19873 23247 19907
rect 23247 19873 23256 19907
rect 23204 19864 23256 19873
rect 23480 19864 23532 19916
rect 26792 19864 26844 19916
rect 24584 19796 24636 19848
rect 25780 19839 25832 19848
rect 25780 19805 25789 19839
rect 25789 19805 25823 19839
rect 25823 19805 25832 19839
rect 25780 19796 25832 19805
rect 12716 19728 12768 19780
rect 13268 19728 13320 19780
rect 14096 19728 14148 19780
rect 11060 19660 11112 19712
rect 13084 19660 13136 19712
rect 15016 19728 15068 19780
rect 20352 19728 20404 19780
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 23572 19660 23624 19712
rect 26700 19660 26752 19712
rect 5536 19558 5588 19610
rect 5600 19558 5652 19610
rect 5664 19558 5716 19610
rect 5728 19558 5780 19610
rect 14644 19558 14696 19610
rect 14708 19558 14760 19610
rect 14772 19558 14824 19610
rect 14836 19558 14888 19610
rect 23752 19558 23804 19610
rect 23816 19558 23868 19610
rect 23880 19558 23932 19610
rect 23944 19558 23996 19610
rect 2320 19456 2372 19508
rect 9956 19456 10008 19508
rect 10692 19456 10744 19508
rect 13728 19456 13780 19508
rect 14464 19456 14516 19508
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 13084 19388 13136 19440
rect 13452 19388 13504 19440
rect 1584 19252 1636 19304
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 5908 19252 5960 19304
rect 6276 19252 6328 19304
rect 6460 19252 6512 19304
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 7380 19295 7432 19304
rect 4804 19184 4856 19236
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 7564 19252 7616 19304
rect 10784 19320 10836 19372
rect 9772 19252 9824 19304
rect 11244 19320 11296 19372
rect 11152 19295 11204 19304
rect 11152 19261 11161 19295
rect 11161 19261 11195 19295
rect 11195 19261 11204 19295
rect 11152 19252 11204 19261
rect 4528 19116 4580 19168
rect 7012 19116 7064 19168
rect 7104 19116 7156 19168
rect 7840 19184 7892 19236
rect 12256 19252 12308 19304
rect 13912 19252 13964 19304
rect 8392 19116 8444 19168
rect 9680 19116 9732 19168
rect 11980 19184 12032 19236
rect 15752 19388 15804 19440
rect 17592 19388 17644 19440
rect 20720 19456 20772 19508
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 15108 19320 15160 19372
rect 22652 19388 22704 19440
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 20352 19320 20404 19372
rect 10876 19116 10928 19168
rect 11060 19116 11112 19168
rect 11612 19116 11664 19168
rect 13360 19116 13412 19168
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15752 19252 15804 19304
rect 18328 19252 18380 19304
rect 18788 19252 18840 19304
rect 20628 19252 20680 19304
rect 20904 19295 20956 19304
rect 20904 19261 20913 19295
rect 20913 19261 20947 19295
rect 20947 19261 20956 19295
rect 20904 19252 20956 19261
rect 14740 19184 14792 19236
rect 14464 19116 14516 19168
rect 17132 19159 17184 19168
rect 17132 19125 17141 19159
rect 17141 19125 17175 19159
rect 17175 19125 17184 19159
rect 17132 19116 17184 19125
rect 20720 19184 20772 19236
rect 23204 19456 23256 19508
rect 21364 19184 21416 19236
rect 22560 19184 22612 19236
rect 25780 19252 25832 19304
rect 26700 19252 26752 19304
rect 27344 19252 27396 19304
rect 23296 19184 23348 19236
rect 23572 19184 23624 19236
rect 22468 19116 22520 19168
rect 22928 19116 22980 19168
rect 23020 19116 23072 19168
rect 24492 19116 24544 19168
rect 24584 19116 24636 19168
rect 10090 19014 10142 19066
rect 10154 19014 10206 19066
rect 10218 19014 10270 19066
rect 10282 19014 10334 19066
rect 19198 19014 19250 19066
rect 19262 19014 19314 19066
rect 19326 19014 19378 19066
rect 19390 19014 19442 19066
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 6276 18912 6328 18964
rect 7380 18912 7432 18964
rect 7472 18912 7524 18964
rect 2872 18844 2924 18896
rect 4528 18887 4580 18896
rect 4528 18853 4537 18887
rect 4537 18853 4571 18887
rect 4571 18853 4580 18887
rect 4528 18844 4580 18853
rect 2320 18776 2372 18828
rect 4252 18819 4304 18828
rect 4252 18785 4261 18819
rect 4261 18785 4295 18819
rect 4295 18785 4304 18819
rect 4252 18776 4304 18785
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 4712 18776 4764 18828
rect 6092 18776 6144 18828
rect 6552 18819 6604 18828
rect 6552 18785 6561 18819
rect 6561 18785 6595 18819
rect 6595 18785 6604 18819
rect 6552 18776 6604 18785
rect 6736 18776 6788 18828
rect 8392 18819 8444 18828
rect 7104 18708 7156 18760
rect 6460 18640 6512 18692
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 2504 18572 2556 18624
rect 6092 18572 6144 18624
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 12348 18844 12400 18896
rect 14096 18912 14148 18964
rect 18236 18912 18288 18964
rect 20076 18912 20128 18964
rect 23296 18955 23348 18964
rect 13268 18844 13320 18896
rect 10232 18776 10284 18828
rect 10324 18776 10376 18828
rect 11888 18819 11940 18828
rect 11888 18785 11897 18819
rect 11897 18785 11931 18819
rect 11931 18785 11940 18819
rect 11888 18776 11940 18785
rect 12992 18819 13044 18828
rect 12992 18785 13001 18819
rect 13001 18785 13035 18819
rect 13035 18785 13044 18819
rect 12992 18776 13044 18785
rect 13360 18819 13412 18828
rect 13360 18785 13369 18819
rect 13369 18785 13403 18819
rect 13403 18785 13412 18819
rect 13360 18776 13412 18785
rect 13912 18776 13964 18828
rect 14740 18819 14792 18828
rect 14740 18785 14749 18819
rect 14749 18785 14783 18819
rect 14783 18785 14792 18819
rect 14740 18776 14792 18785
rect 15016 18776 15068 18828
rect 15936 18819 15988 18828
rect 8392 18640 8444 18692
rect 9956 18640 10008 18692
rect 10416 18640 10468 18692
rect 12256 18708 12308 18760
rect 14464 18708 14516 18760
rect 15108 18751 15160 18760
rect 15108 18717 15117 18751
rect 15117 18717 15151 18751
rect 15151 18717 15160 18751
rect 15108 18708 15160 18717
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 7104 18572 7156 18624
rect 7380 18572 7432 18624
rect 9772 18572 9824 18624
rect 10324 18572 10376 18624
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 13728 18640 13780 18692
rect 17592 18776 17644 18828
rect 17776 18819 17828 18828
rect 17776 18785 17785 18819
rect 17785 18785 17819 18819
rect 17819 18785 17828 18819
rect 17776 18776 17828 18785
rect 23020 18887 23072 18896
rect 17868 18708 17920 18760
rect 18604 18819 18656 18828
rect 18604 18785 18613 18819
rect 18613 18785 18647 18819
rect 18647 18785 18656 18819
rect 18604 18776 18656 18785
rect 20076 18776 20128 18828
rect 20536 18776 20588 18828
rect 20996 18776 21048 18828
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 19800 18708 19852 18760
rect 23020 18853 23029 18887
rect 23029 18853 23063 18887
rect 23063 18853 23072 18887
rect 23020 18844 23072 18853
rect 23296 18921 23305 18955
rect 23305 18921 23339 18955
rect 23339 18921 23348 18955
rect 23296 18912 23348 18921
rect 24768 18912 24820 18964
rect 26240 18912 26292 18964
rect 26792 18955 26844 18964
rect 26792 18921 26801 18955
rect 26801 18921 26835 18955
rect 26835 18921 26844 18955
rect 26792 18912 26844 18921
rect 22928 18819 22980 18828
rect 22928 18785 22937 18819
rect 22937 18785 22971 18819
rect 22971 18785 22980 18819
rect 22928 18776 22980 18785
rect 23204 18776 23256 18828
rect 24400 18776 24452 18828
rect 25320 18844 25372 18896
rect 26976 18844 27028 18896
rect 27528 18887 27580 18896
rect 27528 18853 27537 18887
rect 27537 18853 27571 18887
rect 27571 18853 27580 18887
rect 27528 18844 27580 18853
rect 24492 18708 24544 18760
rect 24768 18708 24820 18760
rect 26240 18819 26292 18828
rect 26240 18785 26249 18819
rect 26249 18785 26283 18819
rect 26283 18785 26292 18819
rect 26240 18776 26292 18785
rect 24124 18640 24176 18692
rect 26608 18819 26660 18828
rect 26608 18785 26617 18819
rect 26617 18785 26651 18819
rect 26651 18785 26660 18819
rect 26608 18776 26660 18785
rect 15200 18572 15252 18624
rect 15384 18615 15436 18624
rect 15384 18581 15393 18615
rect 15393 18581 15427 18615
rect 15427 18581 15436 18615
rect 15384 18572 15436 18581
rect 16580 18572 16632 18624
rect 20260 18572 20312 18624
rect 26240 18572 26292 18624
rect 27620 18615 27672 18624
rect 27620 18581 27629 18615
rect 27629 18581 27663 18615
rect 27663 18581 27672 18615
rect 27620 18572 27672 18581
rect 5536 18470 5588 18522
rect 5600 18470 5652 18522
rect 5664 18470 5716 18522
rect 5728 18470 5780 18522
rect 14644 18470 14696 18522
rect 14708 18470 14760 18522
rect 14772 18470 14824 18522
rect 14836 18470 14888 18522
rect 23752 18470 23804 18522
rect 23816 18470 23868 18522
rect 23880 18470 23932 18522
rect 23944 18470 23996 18522
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 5080 18368 5132 18420
rect 9864 18368 9916 18420
rect 10692 18368 10744 18420
rect 13728 18368 13780 18420
rect 2872 18164 2924 18216
rect 3056 18164 3108 18216
rect 6092 18300 6144 18352
rect 7840 18300 7892 18352
rect 6368 18232 6420 18284
rect 6460 18232 6512 18284
rect 7012 18275 7064 18284
rect 6000 18164 6052 18216
rect 6736 18164 6788 18216
rect 7012 18241 7021 18275
rect 7021 18241 7055 18275
rect 7055 18241 7064 18275
rect 7012 18232 7064 18241
rect 7380 18207 7432 18216
rect 2044 18096 2096 18148
rect 4804 18096 4856 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 4620 18028 4672 18080
rect 6920 18096 6972 18148
rect 7380 18173 7389 18207
rect 7389 18173 7423 18207
rect 7423 18173 7432 18207
rect 7380 18164 7432 18173
rect 7472 18164 7524 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 10876 18164 10928 18216
rect 5908 18071 5960 18080
rect 5908 18037 5917 18071
rect 5917 18037 5951 18071
rect 5951 18037 5960 18071
rect 5908 18028 5960 18037
rect 10508 18096 10560 18148
rect 12992 18300 13044 18352
rect 12256 18207 12308 18216
rect 11612 18096 11664 18148
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 12532 18164 12584 18216
rect 12348 18139 12400 18148
rect 12348 18105 12357 18139
rect 12357 18105 12391 18139
rect 12391 18105 12400 18139
rect 12348 18096 12400 18105
rect 13544 18300 13596 18352
rect 18236 18368 18288 18420
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 20536 18411 20588 18420
rect 20536 18377 20545 18411
rect 20545 18377 20579 18411
rect 20579 18377 20588 18411
rect 20536 18368 20588 18377
rect 20996 18368 21048 18420
rect 24400 18368 24452 18420
rect 27068 18368 27120 18420
rect 15016 18300 15068 18352
rect 15936 18300 15988 18352
rect 18052 18300 18104 18352
rect 13360 18232 13412 18284
rect 14464 18232 14516 18284
rect 18604 18232 18656 18284
rect 15108 18164 15160 18216
rect 15476 18164 15528 18216
rect 13268 18096 13320 18148
rect 13360 18096 13412 18148
rect 13636 18096 13688 18148
rect 16764 18096 16816 18148
rect 18420 18096 18472 18148
rect 19984 18300 20036 18352
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20260 18207 20312 18216
rect 20260 18173 20269 18207
rect 20269 18173 20303 18207
rect 20303 18173 20312 18207
rect 20260 18164 20312 18173
rect 20352 18207 20404 18216
rect 20352 18173 20361 18207
rect 20361 18173 20395 18207
rect 20395 18173 20404 18207
rect 20352 18164 20404 18173
rect 20628 18164 20680 18216
rect 20536 18096 20588 18148
rect 24308 18164 24360 18216
rect 12624 18071 12676 18080
rect 12624 18037 12633 18071
rect 12633 18037 12667 18071
rect 12667 18037 12676 18071
rect 12624 18028 12676 18037
rect 14188 18028 14240 18080
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 16396 18028 16448 18080
rect 17408 18028 17460 18080
rect 21364 18028 21416 18080
rect 22560 18028 22612 18080
rect 25596 18096 25648 18148
rect 25872 18028 25924 18080
rect 27344 18028 27396 18080
rect 10090 17926 10142 17978
rect 10154 17926 10206 17978
rect 10218 17926 10270 17978
rect 10282 17926 10334 17978
rect 19198 17926 19250 17978
rect 19262 17926 19314 17978
rect 19326 17926 19378 17978
rect 19390 17926 19442 17978
rect 3424 17824 3476 17876
rect 4804 17867 4856 17876
rect 4528 17799 4580 17808
rect 4528 17765 4537 17799
rect 4537 17765 4571 17799
rect 4571 17765 4580 17799
rect 4528 17756 4580 17765
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 6920 17824 6972 17876
rect 4068 17688 4120 17740
rect 4344 17688 4396 17740
rect 1400 17620 1452 17672
rect 4712 17688 4764 17740
rect 5908 17756 5960 17808
rect 7564 17824 7616 17876
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 10508 17867 10560 17876
rect 10508 17833 10517 17867
rect 10517 17833 10551 17867
rect 10551 17833 10560 17867
rect 10508 17824 10560 17833
rect 10968 17824 11020 17876
rect 4528 17620 4580 17672
rect 1584 17484 1636 17536
rect 2688 17484 2740 17536
rect 8208 17688 8260 17740
rect 11612 17756 11664 17808
rect 12624 17756 12676 17808
rect 14372 17756 14424 17808
rect 16488 17756 16540 17808
rect 18788 17824 18840 17876
rect 20076 17867 20128 17876
rect 20076 17833 20085 17867
rect 20085 17833 20119 17867
rect 20119 17833 20128 17867
rect 20076 17824 20128 17833
rect 20720 17756 20772 17808
rect 9956 17731 10008 17740
rect 9956 17697 9965 17731
rect 9965 17697 9999 17731
rect 9999 17697 10008 17731
rect 9956 17688 10008 17697
rect 10692 17688 10744 17740
rect 10876 17688 10928 17740
rect 12072 17688 12124 17740
rect 13912 17688 13964 17740
rect 14280 17688 14332 17740
rect 15752 17688 15804 17740
rect 18604 17688 18656 17740
rect 18880 17688 18932 17740
rect 20260 17688 20312 17740
rect 10968 17620 11020 17672
rect 12624 17620 12676 17672
rect 26792 17824 26844 17876
rect 23480 17756 23532 17808
rect 26240 17799 26292 17808
rect 26240 17765 26274 17799
rect 26274 17765 26292 17799
rect 26240 17756 26292 17765
rect 10876 17552 10928 17604
rect 6000 17484 6052 17536
rect 12256 17484 12308 17536
rect 12532 17484 12584 17536
rect 13268 17484 13320 17536
rect 15016 17552 15068 17604
rect 14096 17484 14148 17536
rect 14464 17484 14516 17536
rect 16672 17552 16724 17604
rect 25504 17731 25556 17740
rect 25504 17697 25513 17731
rect 25513 17697 25547 17731
rect 25547 17697 25556 17731
rect 25504 17688 25556 17697
rect 25872 17688 25924 17740
rect 15200 17484 15252 17536
rect 15752 17484 15804 17536
rect 18972 17484 19024 17536
rect 19156 17484 19208 17536
rect 25780 17620 25832 17672
rect 22192 17527 22244 17536
rect 22192 17493 22201 17527
rect 22201 17493 22235 17527
rect 22235 17493 22244 17527
rect 22192 17484 22244 17493
rect 26976 17484 27028 17536
rect 27528 17484 27580 17536
rect 5536 17382 5588 17434
rect 5600 17382 5652 17434
rect 5664 17382 5716 17434
rect 5728 17382 5780 17434
rect 14644 17382 14696 17434
rect 14708 17382 14760 17434
rect 14772 17382 14824 17434
rect 14836 17382 14888 17434
rect 23752 17382 23804 17434
rect 23816 17382 23868 17434
rect 23880 17382 23932 17434
rect 23944 17382 23996 17434
rect 1400 17280 1452 17332
rect 3056 17280 3108 17332
rect 4068 17280 4120 17332
rect 6552 17280 6604 17332
rect 9128 17323 9180 17332
rect 2780 17212 2832 17264
rect 3976 17212 4028 17264
rect 4344 17212 4396 17264
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 10600 17280 10652 17332
rect 12532 17280 12584 17332
rect 25596 17323 25648 17332
rect 7104 17255 7156 17264
rect 7104 17221 7113 17255
rect 7113 17221 7147 17255
rect 7147 17221 7156 17255
rect 7104 17212 7156 17221
rect 16212 17212 16264 17264
rect 19156 17212 19208 17264
rect 2688 17076 2740 17128
rect 3608 17119 3660 17128
rect 3148 17008 3200 17060
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 3976 17119 4028 17128
rect 3976 17085 3985 17119
rect 3985 17085 4019 17119
rect 4019 17085 4028 17119
rect 3976 17076 4028 17085
rect 4344 17008 4396 17060
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 4620 17076 4672 17085
rect 8852 17144 8904 17196
rect 7380 17076 7432 17128
rect 8024 17076 8076 17128
rect 2964 16940 3016 16992
rect 4620 16940 4672 16992
rect 7472 17008 7524 17060
rect 7840 17008 7892 17060
rect 9036 17051 9088 17060
rect 9036 17017 9045 17051
rect 9045 17017 9079 17051
rect 9079 17017 9088 17051
rect 9036 17008 9088 17017
rect 9680 17008 9732 17060
rect 9864 16940 9916 16992
rect 12348 17144 12400 17196
rect 11888 17076 11940 17128
rect 17408 17144 17460 17196
rect 17684 17144 17736 17196
rect 17776 17144 17828 17196
rect 25596 17289 25605 17323
rect 25605 17289 25639 17323
rect 25639 17289 25648 17323
rect 25596 17280 25648 17289
rect 20720 17212 20772 17264
rect 26884 17255 26936 17264
rect 19616 17144 19668 17196
rect 11520 17008 11572 17060
rect 13544 16940 13596 16992
rect 13636 16940 13688 16992
rect 14188 17008 14240 17060
rect 20260 17076 20312 17128
rect 22192 17144 22244 17196
rect 15476 17008 15528 17060
rect 16304 17008 16356 17060
rect 18236 17008 18288 17060
rect 21456 17076 21508 17128
rect 21548 17076 21600 17128
rect 23940 17076 23992 17128
rect 26884 17221 26893 17255
rect 26893 17221 26927 17255
rect 26927 17221 26936 17255
rect 26884 17212 26936 17221
rect 25320 17119 25372 17128
rect 21088 17008 21140 17060
rect 22744 17051 22796 17060
rect 22744 17017 22753 17051
rect 22753 17017 22787 17051
rect 22787 17017 22796 17051
rect 22744 17008 22796 17017
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 27344 17144 27396 17196
rect 26700 17119 26752 17128
rect 26700 17085 26709 17119
rect 26709 17085 26743 17119
rect 26743 17085 26752 17119
rect 26700 17076 26752 17085
rect 15752 16940 15804 16992
rect 16488 16940 16540 16992
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 17408 16940 17460 16992
rect 17960 16940 18012 16992
rect 18052 16940 18104 16992
rect 20720 16940 20772 16992
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 22468 16940 22520 16992
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 24952 16940 25004 16992
rect 25504 16940 25556 16992
rect 10090 16838 10142 16890
rect 10154 16838 10206 16890
rect 10218 16838 10270 16890
rect 10282 16838 10334 16890
rect 19198 16838 19250 16890
rect 19262 16838 19314 16890
rect 19326 16838 19378 16890
rect 19390 16838 19442 16890
rect 1768 16736 1820 16788
rect 2412 16736 2464 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 3608 16736 3660 16788
rect 6276 16736 6328 16788
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 2964 16668 3016 16720
rect 4436 16668 4488 16720
rect 5356 16668 5408 16720
rect 6000 16668 6052 16720
rect 6460 16668 6512 16720
rect 6644 16668 6696 16720
rect 10600 16736 10652 16788
rect 10876 16779 10928 16788
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 10968 16736 11020 16788
rect 12348 16736 12400 16788
rect 15476 16736 15528 16788
rect 2780 16532 2832 16584
rect 3148 16600 3200 16652
rect 3884 16600 3936 16652
rect 7012 16600 7064 16652
rect 12072 16668 12124 16720
rect 12624 16711 12676 16720
rect 12624 16677 12633 16711
rect 12633 16677 12667 16711
rect 12667 16677 12676 16711
rect 12624 16668 12676 16677
rect 13452 16668 13504 16720
rect 16488 16736 16540 16788
rect 17960 16736 18012 16788
rect 18052 16736 18104 16788
rect 19708 16736 19760 16788
rect 21456 16736 21508 16788
rect 23940 16779 23992 16788
rect 23940 16745 23949 16779
rect 23949 16745 23983 16779
rect 23983 16745 23992 16779
rect 23940 16736 23992 16745
rect 24492 16736 24544 16788
rect 25872 16736 25924 16788
rect 26148 16736 26200 16788
rect 17316 16668 17368 16720
rect 9772 16643 9824 16652
rect 9772 16609 9806 16643
rect 9806 16609 9824 16643
rect 1860 16396 1912 16448
rect 7104 16464 7156 16516
rect 9772 16600 9824 16609
rect 11520 16600 11572 16652
rect 12532 16600 12584 16652
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 13544 16600 13596 16652
rect 14464 16600 14516 16652
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 18788 16668 18840 16720
rect 20904 16668 20956 16720
rect 23112 16668 23164 16720
rect 26608 16668 26660 16720
rect 15752 16600 15804 16609
rect 17868 16643 17920 16652
rect 17868 16609 17902 16643
rect 17902 16609 17920 16643
rect 17868 16600 17920 16609
rect 19800 16600 19852 16652
rect 15016 16532 15068 16584
rect 12716 16396 12768 16448
rect 20076 16396 20128 16448
rect 20260 16600 20312 16652
rect 22468 16600 22520 16652
rect 25596 16643 25648 16652
rect 25596 16609 25605 16643
rect 25605 16609 25639 16643
rect 25639 16609 25648 16643
rect 25596 16600 25648 16609
rect 25780 16600 25832 16652
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 24584 16396 24636 16448
rect 5536 16294 5588 16346
rect 5600 16294 5652 16346
rect 5664 16294 5716 16346
rect 5728 16294 5780 16346
rect 14644 16294 14696 16346
rect 14708 16294 14760 16346
rect 14772 16294 14824 16346
rect 14836 16294 14888 16346
rect 23752 16294 23804 16346
rect 23816 16294 23868 16346
rect 23880 16294 23932 16346
rect 23944 16294 23996 16346
rect 2136 16192 2188 16244
rect 15200 16192 15252 16244
rect 18604 16192 18656 16244
rect 20628 16192 20680 16244
rect 21088 16192 21140 16244
rect 21272 16192 21324 16244
rect 24768 16192 24820 16244
rect 25228 16192 25280 16244
rect 26516 16192 26568 16244
rect 6368 16124 6420 16176
rect 6460 16124 6512 16176
rect 13452 16167 13504 16176
rect 2044 15988 2096 16040
rect 2228 15988 2280 16040
rect 3792 16031 3844 16040
rect 3792 15997 3801 16031
rect 3801 15997 3835 16031
rect 3835 15997 3844 16031
rect 3792 15988 3844 15997
rect 6092 16056 6144 16108
rect 4344 15920 4396 15972
rect 5816 15988 5868 16040
rect 4160 15895 4212 15904
rect 4160 15861 4169 15895
rect 4169 15861 4203 15895
rect 4203 15861 4212 15895
rect 4160 15852 4212 15861
rect 4896 15963 4948 15972
rect 4896 15929 4905 15963
rect 4905 15929 4939 15963
rect 4939 15929 4948 15963
rect 4896 15920 4948 15929
rect 5908 15920 5960 15972
rect 6736 16056 6788 16108
rect 13452 16133 13461 16167
rect 13461 16133 13495 16167
rect 13495 16133 13504 16167
rect 13452 16124 13504 16133
rect 15936 16167 15988 16176
rect 15936 16133 15945 16167
rect 15945 16133 15979 16167
rect 15979 16133 15988 16167
rect 15936 16124 15988 16133
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 7104 15988 7156 15997
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 12716 15988 12768 16040
rect 6644 15920 6696 15972
rect 4988 15852 5040 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5356 15852 5408 15904
rect 7840 15920 7892 15972
rect 8576 15920 8628 15972
rect 7104 15852 7156 15904
rect 9864 15895 9916 15904
rect 9864 15861 9873 15895
rect 9873 15861 9907 15895
rect 9907 15861 9916 15895
rect 13452 15988 13504 16040
rect 17868 16167 17920 16176
rect 17868 16133 17877 16167
rect 17877 16133 17911 16167
rect 17911 16133 17920 16167
rect 17868 16124 17920 16133
rect 18236 16124 18288 16176
rect 23388 16124 23440 16176
rect 24584 16099 24636 16108
rect 16304 15988 16356 16040
rect 17868 15988 17920 16040
rect 18604 15988 18656 16040
rect 18972 15988 19024 16040
rect 15016 15920 15068 15972
rect 17408 15920 17460 15972
rect 18052 15920 18104 15972
rect 18328 15920 18380 15972
rect 19616 16031 19668 16040
rect 19616 15997 19625 16031
rect 19625 15997 19659 16031
rect 19659 15997 19668 16031
rect 19616 15988 19668 15997
rect 20444 15988 20496 16040
rect 23480 15988 23532 16040
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 25320 15988 25372 16040
rect 19708 15920 19760 15972
rect 20904 15920 20956 15972
rect 20996 15920 21048 15972
rect 21916 15920 21968 15972
rect 23572 15963 23624 15972
rect 23572 15929 23581 15963
rect 23581 15929 23615 15963
rect 23615 15929 23624 15963
rect 23572 15920 23624 15929
rect 24860 15963 24912 15972
rect 24860 15929 24894 15963
rect 24894 15929 24912 15963
rect 24860 15920 24912 15929
rect 26884 15920 26936 15972
rect 9864 15852 9916 15861
rect 13728 15852 13780 15904
rect 20812 15852 20864 15904
rect 22284 15852 22336 15904
rect 10090 15750 10142 15802
rect 10154 15750 10206 15802
rect 10218 15750 10270 15802
rect 10282 15750 10334 15802
rect 19198 15750 19250 15802
rect 19262 15750 19314 15802
rect 19326 15750 19378 15802
rect 19390 15750 19442 15802
rect 2320 15648 2372 15700
rect 6000 15648 6052 15700
rect 6276 15648 6328 15700
rect 5172 15580 5224 15632
rect 6736 15580 6788 15632
rect 7288 15580 7340 15632
rect 7656 15580 7708 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 6460 15512 6512 15564
rect 6920 15512 6972 15564
rect 9772 15648 9824 15700
rect 10692 15648 10744 15700
rect 12900 15580 12952 15632
rect 10876 15555 10928 15564
rect 5816 15376 5868 15428
rect 10692 15444 10744 15496
rect 10876 15521 10902 15555
rect 10902 15521 10928 15555
rect 10876 15512 10928 15521
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 14372 15580 14424 15632
rect 16488 15580 16540 15632
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 15292 15512 15344 15564
rect 17040 15512 17092 15564
rect 10968 15444 11020 15496
rect 12072 15444 12124 15496
rect 17960 15512 18012 15564
rect 20076 15580 20128 15632
rect 21916 15623 21968 15632
rect 20260 15555 20312 15564
rect 20260 15521 20294 15555
rect 20294 15521 20312 15555
rect 21916 15589 21925 15623
rect 21925 15589 21959 15623
rect 21959 15589 21968 15623
rect 21916 15580 21968 15589
rect 23388 15648 23440 15700
rect 26516 15648 26568 15700
rect 27252 15648 27304 15700
rect 25596 15580 25648 15632
rect 20260 15512 20312 15521
rect 2320 15308 2372 15360
rect 4896 15308 4948 15360
rect 6184 15308 6236 15360
rect 9036 15376 9088 15428
rect 10876 15376 10928 15428
rect 11060 15419 11112 15428
rect 11060 15385 11069 15419
rect 11069 15385 11103 15419
rect 11103 15385 11112 15419
rect 11060 15376 11112 15385
rect 14188 15376 14240 15428
rect 12808 15308 12860 15360
rect 13176 15351 13228 15360
rect 13176 15317 13185 15351
rect 13185 15317 13219 15351
rect 13219 15317 13228 15351
rect 13176 15308 13228 15317
rect 13820 15308 13872 15360
rect 15752 15376 15804 15428
rect 17224 15376 17276 15428
rect 17868 15376 17920 15428
rect 17408 15308 17460 15360
rect 18052 15308 18104 15360
rect 18880 15351 18932 15360
rect 18880 15317 18889 15351
rect 18889 15317 18923 15351
rect 18923 15317 18932 15351
rect 18880 15308 18932 15317
rect 23388 15512 23440 15564
rect 24952 15512 25004 15564
rect 27068 15555 27120 15564
rect 27068 15521 27077 15555
rect 27077 15521 27111 15555
rect 27111 15521 27120 15555
rect 27068 15512 27120 15521
rect 27252 15555 27304 15564
rect 27252 15521 27261 15555
rect 27261 15521 27295 15555
rect 27295 15521 27304 15555
rect 27252 15512 27304 15521
rect 27436 15555 27488 15564
rect 27436 15521 27445 15555
rect 27445 15521 27479 15555
rect 27479 15521 27488 15555
rect 27436 15512 27488 15521
rect 22100 15419 22152 15428
rect 22100 15385 22109 15419
rect 22109 15385 22143 15419
rect 22143 15385 22152 15419
rect 22100 15376 22152 15385
rect 20720 15308 20772 15360
rect 21916 15308 21968 15360
rect 25412 15308 25464 15360
rect 26700 15308 26752 15360
rect 5536 15206 5588 15258
rect 5600 15206 5652 15258
rect 5664 15206 5716 15258
rect 5728 15206 5780 15258
rect 14644 15206 14696 15258
rect 14708 15206 14760 15258
rect 14772 15206 14824 15258
rect 14836 15206 14888 15258
rect 23752 15206 23804 15258
rect 23816 15206 23868 15258
rect 23880 15206 23932 15258
rect 23944 15206 23996 15258
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 7104 15104 7156 15156
rect 13084 15104 13136 15156
rect 13360 15104 13412 15156
rect 14464 15104 14516 15156
rect 23204 15104 23256 15156
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 23388 15104 23440 15113
rect 24860 15104 24912 15156
rect 27436 15104 27488 15156
rect 9220 15036 9272 15088
rect 6920 14968 6972 15020
rect 9128 14968 9180 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 2780 14900 2832 14952
rect 4160 14900 4212 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 8760 14943 8812 14952
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 9312 14943 9364 14952
rect 8944 14832 8996 14884
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 9496 15036 9548 15088
rect 10692 15079 10744 15088
rect 10692 15045 10701 15079
rect 10701 15045 10735 15079
rect 10735 15045 10744 15079
rect 10692 15036 10744 15045
rect 15292 15079 15344 15088
rect 15292 15045 15301 15079
rect 15301 15045 15335 15079
rect 15335 15045 15344 15079
rect 15292 15036 15344 15045
rect 18512 15036 18564 15088
rect 20260 15079 20312 15088
rect 11336 14968 11388 15020
rect 11520 14968 11572 15020
rect 14096 14968 14148 15020
rect 9680 14900 9732 14952
rect 10416 14832 10468 14884
rect 11428 14832 11480 14884
rect 12624 14900 12676 14952
rect 14188 14900 14240 14952
rect 14740 14943 14792 14952
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 14924 14900 14976 14909
rect 17316 14968 17368 15020
rect 17960 14968 18012 15020
rect 15292 14900 15344 14952
rect 7472 14764 7524 14816
rect 7932 14764 7984 14816
rect 14832 14832 14884 14884
rect 15752 14832 15804 14884
rect 17592 14943 17644 14952
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 18788 14968 18840 15020
rect 18328 14900 18380 14952
rect 14464 14764 14516 14816
rect 14740 14764 14792 14816
rect 16856 14764 16908 14816
rect 18880 14832 18932 14884
rect 20260 15045 20269 15079
rect 20269 15045 20303 15079
rect 20303 15045 20312 15079
rect 20260 15036 20312 15045
rect 21640 15079 21692 15088
rect 21640 15045 21649 15079
rect 21649 15045 21683 15079
rect 21683 15045 21692 15079
rect 21640 15036 21692 15045
rect 22100 15036 22152 15088
rect 19524 14900 19576 14952
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 18328 14764 18380 14816
rect 19708 14764 19760 14816
rect 19984 14875 20036 14884
rect 19984 14841 19993 14875
rect 19993 14841 20027 14875
rect 20027 14841 20036 14875
rect 21088 14943 21140 14952
rect 21088 14909 21097 14943
rect 21097 14909 21131 14943
rect 21131 14909 21140 14943
rect 21088 14900 21140 14909
rect 21272 14943 21324 14952
rect 21272 14909 21281 14943
rect 21281 14909 21315 14943
rect 21315 14909 21324 14943
rect 21272 14900 21324 14909
rect 21364 14875 21416 14884
rect 19984 14832 20036 14841
rect 21364 14841 21373 14875
rect 21373 14841 21407 14875
rect 21407 14841 21416 14875
rect 21364 14832 21416 14841
rect 22928 14900 22980 14952
rect 23480 15036 23532 15088
rect 23296 14900 23348 14952
rect 23480 14900 23532 14952
rect 23572 14832 23624 14884
rect 24216 14943 24268 14952
rect 24216 14909 24225 14943
rect 24225 14909 24259 14943
rect 24259 14909 24268 14943
rect 24216 14900 24268 14909
rect 25228 14900 25280 14952
rect 24584 14832 24636 14884
rect 25136 14832 25188 14884
rect 25412 14832 25464 14884
rect 26700 14900 26752 14952
rect 26056 14832 26108 14884
rect 22468 14764 22520 14816
rect 10090 14662 10142 14714
rect 10154 14662 10206 14714
rect 10218 14662 10270 14714
rect 10282 14662 10334 14714
rect 19198 14662 19250 14714
rect 19262 14662 19314 14714
rect 19326 14662 19378 14714
rect 19390 14662 19442 14714
rect 7104 14560 7156 14612
rect 2412 14492 2464 14544
rect 8392 14560 8444 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 8668 14560 8720 14612
rect 9404 14560 9456 14612
rect 9864 14560 9916 14612
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 4344 14424 4396 14476
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 1952 14356 2004 14408
rect 7656 14424 7708 14476
rect 7840 14356 7892 14408
rect 9680 14424 9732 14476
rect 11060 14560 11112 14612
rect 10876 14492 10928 14544
rect 10416 14467 10468 14476
rect 10416 14433 10425 14467
rect 10425 14433 10459 14467
rect 10459 14433 10468 14467
rect 10416 14424 10468 14433
rect 10968 14424 11020 14476
rect 11152 14424 11204 14476
rect 2044 14331 2096 14340
rect 2044 14297 2053 14331
rect 2053 14297 2087 14331
rect 2087 14297 2096 14331
rect 2044 14288 2096 14297
rect 6736 14288 6788 14340
rect 5080 14220 5132 14272
rect 5356 14220 5408 14272
rect 7656 14220 7708 14272
rect 9128 14356 9180 14408
rect 10784 14356 10836 14408
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 8576 14288 8628 14340
rect 22284 14560 22336 14612
rect 22468 14560 22520 14612
rect 15016 14535 15068 14544
rect 15016 14501 15025 14535
rect 15025 14501 15059 14535
rect 15059 14501 15068 14535
rect 15016 14492 15068 14501
rect 15936 14492 15988 14544
rect 16304 14492 16356 14544
rect 16764 14492 16816 14544
rect 13452 14424 13504 14476
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 14924 14467 14976 14476
rect 14464 14356 14516 14408
rect 14924 14433 14933 14467
rect 14933 14433 14967 14467
rect 14967 14433 14976 14467
rect 14924 14424 14976 14433
rect 15292 14424 15344 14476
rect 15660 14424 15712 14476
rect 16120 14424 16172 14476
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 18328 14492 18380 14544
rect 19616 14492 19668 14544
rect 21640 14492 21692 14544
rect 25596 14535 25648 14544
rect 25596 14501 25605 14535
rect 25605 14501 25639 14535
rect 25639 14501 25648 14535
rect 25596 14492 25648 14501
rect 17224 14467 17276 14476
rect 17224 14433 17233 14467
rect 17233 14433 17267 14467
rect 17267 14433 17276 14467
rect 17408 14467 17460 14476
rect 17224 14424 17276 14433
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 18052 14424 18104 14476
rect 18512 14424 18564 14476
rect 20628 14424 20680 14476
rect 20720 14424 20772 14476
rect 21824 14424 21876 14476
rect 23204 14424 23256 14476
rect 25504 14467 25556 14476
rect 25504 14433 25513 14467
rect 25513 14433 25547 14467
rect 25547 14433 25556 14467
rect 25504 14424 25556 14433
rect 27436 14424 27488 14476
rect 18880 14356 18932 14408
rect 18972 14356 19024 14408
rect 20812 14356 20864 14408
rect 8668 14220 8720 14272
rect 8944 14220 8996 14272
rect 9956 14220 10008 14272
rect 10416 14220 10468 14272
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 13452 14288 13504 14340
rect 12992 14220 13044 14272
rect 13728 14263 13780 14272
rect 13728 14229 13737 14263
rect 13737 14229 13771 14263
rect 13771 14229 13780 14263
rect 13728 14220 13780 14229
rect 15200 14220 15252 14272
rect 17500 14220 17552 14272
rect 18052 14220 18104 14272
rect 20536 14288 20588 14340
rect 23112 14288 23164 14340
rect 25780 14220 25832 14272
rect 26056 14288 26108 14340
rect 27068 14220 27120 14272
rect 5536 14118 5588 14170
rect 5600 14118 5652 14170
rect 5664 14118 5716 14170
rect 5728 14118 5780 14170
rect 14644 14118 14696 14170
rect 14708 14118 14760 14170
rect 14772 14118 14824 14170
rect 14836 14118 14888 14170
rect 23752 14118 23804 14170
rect 23816 14118 23868 14170
rect 23880 14118 23932 14170
rect 23944 14118 23996 14170
rect 7104 14016 7156 14068
rect 8484 14016 8536 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 11336 14016 11388 14068
rect 23112 14016 23164 14068
rect 23204 14016 23256 14068
rect 24952 14059 25004 14068
rect 4344 13948 4396 14000
rect 5356 13948 5408 14000
rect 5540 13948 5592 14000
rect 6644 13948 6696 14000
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 3240 13880 3292 13932
rect 2412 13812 2464 13864
rect 4988 13880 5040 13932
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 5908 13880 5960 13932
rect 2228 13787 2280 13796
rect 2228 13753 2237 13787
rect 2237 13753 2271 13787
rect 2271 13753 2280 13787
rect 2228 13744 2280 13753
rect 4252 13744 4304 13796
rect 6828 13744 6880 13796
rect 6920 13787 6972 13796
rect 6920 13753 6929 13787
rect 6929 13753 6963 13787
rect 6963 13753 6972 13787
rect 7656 13812 7708 13864
rect 10324 13812 10376 13864
rect 11060 13948 11112 14000
rect 13452 13991 13504 14000
rect 13452 13957 13461 13991
rect 13461 13957 13495 13991
rect 13495 13957 13504 13991
rect 13452 13948 13504 13957
rect 14188 13948 14240 14000
rect 13084 13880 13136 13932
rect 16028 13923 16080 13932
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 10968 13855 11020 13864
rect 10968 13821 10977 13855
rect 10977 13821 11011 13855
rect 11011 13821 11020 13855
rect 10968 13812 11020 13821
rect 11336 13812 11388 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 12164 13812 12216 13864
rect 13912 13812 13964 13864
rect 14372 13812 14424 13864
rect 16028 13889 16037 13923
rect 16037 13889 16071 13923
rect 16071 13889 16080 13923
rect 16028 13880 16080 13889
rect 19708 13880 19760 13932
rect 20076 13880 20128 13932
rect 15108 13855 15160 13864
rect 15108 13821 15141 13855
rect 15141 13821 15160 13855
rect 15108 13812 15160 13821
rect 17040 13812 17092 13864
rect 18880 13812 18932 13864
rect 20260 13855 20312 13864
rect 20260 13821 20269 13855
rect 20269 13821 20303 13855
rect 20303 13821 20312 13855
rect 20260 13812 20312 13821
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 20904 13812 20956 13864
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 25688 14016 25740 14068
rect 26056 14016 26108 14068
rect 25412 13948 25464 14000
rect 26148 13991 26200 14000
rect 26148 13957 26157 13991
rect 26157 13957 26191 13991
rect 26191 13957 26200 13991
rect 26148 13948 26200 13957
rect 6920 13744 6972 13753
rect 10692 13744 10744 13796
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 6000 13676 6052 13728
rect 11520 13744 11572 13796
rect 14280 13744 14332 13796
rect 14464 13744 14516 13796
rect 12992 13676 13044 13728
rect 15568 13744 15620 13796
rect 16488 13744 16540 13796
rect 17960 13744 18012 13796
rect 18328 13744 18380 13796
rect 20996 13744 21048 13796
rect 24308 13812 24360 13864
rect 24584 13855 24636 13864
rect 24584 13821 24593 13855
rect 24593 13821 24627 13855
rect 24627 13821 24636 13855
rect 24584 13812 24636 13821
rect 26516 13880 26568 13932
rect 25780 13812 25832 13864
rect 23664 13787 23716 13796
rect 23664 13753 23673 13787
rect 23673 13753 23707 13787
rect 23707 13753 23716 13787
rect 23664 13744 23716 13753
rect 15108 13676 15160 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 19064 13676 19116 13728
rect 20904 13676 20956 13728
rect 23388 13676 23440 13728
rect 10090 13574 10142 13626
rect 10154 13574 10206 13626
rect 10218 13574 10270 13626
rect 10282 13574 10334 13626
rect 19198 13574 19250 13626
rect 19262 13574 19314 13626
rect 19326 13574 19378 13626
rect 19390 13574 19442 13626
rect 2228 13472 2280 13524
rect 2504 13404 2556 13456
rect 4160 13472 4212 13524
rect 5080 13472 5132 13524
rect 6828 13472 6880 13524
rect 8300 13472 8352 13524
rect 9312 13472 9364 13524
rect 10600 13472 10652 13524
rect 12624 13515 12676 13524
rect 5908 13404 5960 13456
rect 9588 13447 9640 13456
rect 5080 13336 5132 13388
rect 7472 13379 7524 13388
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 7656 13336 7708 13388
rect 8300 13379 8352 13388
rect 6920 13268 6972 13320
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 9588 13413 9597 13447
rect 9597 13413 9631 13447
rect 9631 13413 9640 13447
rect 9588 13404 9640 13413
rect 9772 13336 9824 13388
rect 10416 13379 10468 13388
rect 10416 13345 10425 13379
rect 10425 13345 10459 13379
rect 10459 13345 10468 13379
rect 10416 13336 10468 13345
rect 10600 13379 10652 13388
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 12624 13481 12633 13515
rect 12633 13481 12667 13515
rect 12667 13481 12676 13515
rect 12624 13472 12676 13481
rect 15108 13472 15160 13524
rect 15200 13404 15252 13456
rect 15936 13472 15988 13524
rect 16304 13404 16356 13456
rect 17960 13472 18012 13524
rect 18972 13472 19024 13524
rect 17040 13336 17092 13388
rect 19064 13404 19116 13456
rect 21088 13447 21140 13456
rect 21088 13413 21097 13447
rect 21097 13413 21131 13447
rect 21131 13413 21140 13447
rect 21088 13404 21140 13413
rect 18236 13379 18288 13388
rect 10692 13268 10744 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 17316 13268 17368 13320
rect 18236 13345 18245 13379
rect 18245 13345 18279 13379
rect 18279 13345 18288 13379
rect 18236 13336 18288 13345
rect 18880 13379 18932 13388
rect 18880 13345 18889 13379
rect 18889 13345 18923 13379
rect 18923 13345 18932 13379
rect 18880 13336 18932 13345
rect 18604 13268 18656 13320
rect 21088 13268 21140 13320
rect 2780 13132 2832 13184
rect 5080 13132 5132 13184
rect 7288 13200 7340 13252
rect 7472 13200 7524 13252
rect 9036 13200 9088 13252
rect 10416 13200 10468 13252
rect 10784 13200 10836 13252
rect 6644 13132 6696 13184
rect 7656 13132 7708 13184
rect 10968 13132 11020 13184
rect 18052 13200 18104 13252
rect 18972 13243 19024 13252
rect 11612 13132 11664 13184
rect 13728 13132 13780 13184
rect 15936 13132 15988 13184
rect 16672 13132 16724 13184
rect 17684 13132 17736 13184
rect 18420 13132 18472 13184
rect 18972 13209 18981 13243
rect 18981 13209 19015 13243
rect 19015 13209 19024 13243
rect 18972 13200 19024 13209
rect 20812 13200 20864 13252
rect 22100 13336 22152 13388
rect 23296 13336 23348 13388
rect 24308 13472 24360 13524
rect 25228 13472 25280 13524
rect 25412 13404 25464 13456
rect 22560 13268 22612 13320
rect 24124 13336 24176 13388
rect 24860 13336 24912 13388
rect 26976 13336 27028 13388
rect 25136 13268 25188 13320
rect 24216 13200 24268 13252
rect 23480 13132 23532 13184
rect 5536 13030 5588 13082
rect 5600 13030 5652 13082
rect 5664 13030 5716 13082
rect 5728 13030 5780 13082
rect 14644 13030 14696 13082
rect 14708 13030 14760 13082
rect 14772 13030 14824 13082
rect 14836 13030 14888 13082
rect 23752 13030 23804 13082
rect 23816 13030 23868 13082
rect 23880 13030 23932 13082
rect 23944 13030 23996 13082
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 2780 12792 2832 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 4068 12724 4120 12776
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 5448 12724 5500 12776
rect 8300 12928 8352 12980
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 5724 12860 5776 12912
rect 6552 12860 6604 12912
rect 6644 12792 6696 12844
rect 5908 12724 5960 12776
rect 6368 12724 6420 12776
rect 8484 12724 8536 12776
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 10416 12860 10468 12912
rect 10600 12860 10652 12912
rect 10968 12903 11020 12912
rect 10968 12869 10977 12903
rect 10977 12869 11011 12903
rect 11011 12869 11020 12903
rect 10968 12860 11020 12869
rect 11336 12928 11388 12980
rect 13912 12928 13964 12980
rect 14096 12928 14148 12980
rect 11704 12860 11756 12912
rect 12072 12860 12124 12912
rect 12256 12860 12308 12912
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 5724 12588 5776 12640
rect 7196 12656 7248 12708
rect 7840 12656 7892 12708
rect 6092 12588 6144 12640
rect 6644 12588 6696 12640
rect 6736 12588 6788 12640
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 13544 12860 13596 12912
rect 15568 12928 15620 12980
rect 18880 12928 18932 12980
rect 9864 12724 9916 12733
rect 10876 12724 10928 12776
rect 13452 12724 13504 12776
rect 14280 12724 14332 12776
rect 14464 12724 14516 12776
rect 14188 12656 14240 12708
rect 9680 12588 9732 12640
rect 14096 12588 14148 12640
rect 16488 12792 16540 12844
rect 17408 12792 17460 12844
rect 17684 12860 17736 12912
rect 20260 12860 20312 12912
rect 21916 12792 21968 12844
rect 15292 12724 15344 12776
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 14924 12656 14976 12708
rect 17592 12767 17644 12776
rect 17592 12733 17601 12767
rect 17601 12733 17635 12767
rect 17635 12733 17644 12767
rect 17592 12724 17644 12733
rect 18236 12724 18288 12776
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 19616 12767 19668 12776
rect 18328 12724 18380 12733
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 19708 12724 19760 12776
rect 24952 12724 25004 12776
rect 25136 12767 25188 12776
rect 25136 12733 25145 12767
rect 25145 12733 25179 12767
rect 25179 12733 25188 12767
rect 25136 12724 25188 12733
rect 19800 12699 19852 12708
rect 19800 12665 19809 12699
rect 19809 12665 19843 12699
rect 19843 12665 19852 12699
rect 19800 12656 19852 12665
rect 20996 12656 21048 12708
rect 23664 12656 23716 12708
rect 25780 12656 25832 12708
rect 16672 12588 16724 12640
rect 16764 12588 16816 12640
rect 17408 12588 17460 12640
rect 20352 12588 20404 12640
rect 20628 12588 20680 12640
rect 21640 12631 21692 12640
rect 21640 12597 21649 12631
rect 21649 12597 21683 12631
rect 21683 12597 21692 12631
rect 21640 12588 21692 12597
rect 24400 12631 24452 12640
rect 24400 12597 24409 12631
rect 24409 12597 24443 12631
rect 24443 12597 24452 12631
rect 24400 12588 24452 12597
rect 25504 12588 25556 12640
rect 10090 12486 10142 12538
rect 10154 12486 10206 12538
rect 10218 12486 10270 12538
rect 10282 12486 10334 12538
rect 19198 12486 19250 12538
rect 19262 12486 19314 12538
rect 19326 12486 19378 12538
rect 19390 12486 19442 12538
rect 2688 12316 2740 12368
rect 3700 12248 3752 12300
rect 3976 12248 4028 12300
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 4896 12291 4948 12300
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 8024 12384 8076 12436
rect 8576 12316 8628 12368
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 10692 12384 10744 12436
rect 11704 12427 11756 12436
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 11980 12384 12032 12436
rect 14004 12384 14056 12436
rect 14924 12427 14976 12436
rect 14924 12393 14933 12427
rect 14933 12393 14967 12427
rect 14967 12393 14976 12427
rect 14924 12384 14976 12393
rect 16212 12384 16264 12436
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 11336 12316 11388 12368
rect 13820 12316 13872 12368
rect 14188 12316 14240 12368
rect 10692 12248 10744 12300
rect 12992 12291 13044 12300
rect 3424 12044 3476 12096
rect 7380 12180 7432 12232
rect 10784 12180 10836 12232
rect 10876 12180 10928 12232
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 15016 12248 15068 12300
rect 15844 12316 15896 12368
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 16028 12291 16080 12300
rect 15752 12248 15804 12257
rect 16028 12257 16037 12291
rect 16037 12257 16071 12291
rect 16071 12257 16080 12291
rect 16028 12248 16080 12257
rect 16580 12248 16632 12300
rect 17316 12384 17368 12436
rect 18236 12384 18288 12436
rect 19800 12384 19852 12436
rect 16948 12316 17000 12368
rect 6276 12112 6328 12164
rect 4988 12044 5040 12096
rect 12072 12112 12124 12164
rect 12716 12112 12768 12164
rect 15844 12112 15896 12164
rect 16856 12112 16908 12164
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 10324 12044 10376 12053
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 12256 12087 12308 12096
rect 12256 12053 12265 12087
rect 12265 12053 12299 12087
rect 12299 12053 12308 12087
rect 12256 12044 12308 12053
rect 13360 12044 13412 12096
rect 16580 12044 16632 12096
rect 17040 12044 17092 12096
rect 17592 12316 17644 12368
rect 21272 12316 21324 12368
rect 22100 12384 22152 12436
rect 22560 12427 22612 12436
rect 22560 12393 22569 12427
rect 22569 12393 22603 12427
rect 22603 12393 22612 12427
rect 22560 12384 22612 12393
rect 23480 12384 23532 12436
rect 23664 12427 23716 12436
rect 23664 12393 23673 12427
rect 23673 12393 23707 12427
rect 23707 12393 23716 12427
rect 23664 12384 23716 12393
rect 24216 12427 24268 12436
rect 24216 12393 24225 12427
rect 24225 12393 24259 12427
rect 24259 12393 24268 12427
rect 24216 12384 24268 12393
rect 25780 12427 25832 12436
rect 25780 12393 25789 12427
rect 25789 12393 25823 12427
rect 25823 12393 25832 12427
rect 25780 12384 25832 12393
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 19064 12248 19116 12300
rect 20720 12248 20772 12300
rect 21180 12248 21232 12300
rect 21456 12248 21508 12300
rect 21640 12248 21692 12300
rect 24768 12316 24820 12368
rect 26332 12316 26384 12368
rect 26976 12316 27028 12368
rect 17592 12180 17644 12232
rect 19616 12180 19668 12232
rect 22652 12180 22704 12232
rect 24400 12248 24452 12300
rect 25320 12248 25372 12300
rect 25504 12291 25556 12300
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 27712 12291 27764 12300
rect 24216 12180 24268 12232
rect 27712 12257 27721 12291
rect 27721 12257 27755 12291
rect 27755 12257 27764 12291
rect 27712 12248 27764 12257
rect 18696 12112 18748 12164
rect 23572 12112 23624 12164
rect 24768 12112 24820 12164
rect 18144 12044 18196 12096
rect 25320 12044 25372 12096
rect 26884 12087 26936 12096
rect 26884 12053 26893 12087
rect 26893 12053 26927 12087
rect 26927 12053 26936 12087
rect 26884 12044 26936 12053
rect 5536 11942 5588 11994
rect 5600 11942 5652 11994
rect 5664 11942 5716 11994
rect 5728 11942 5780 11994
rect 14644 11942 14696 11994
rect 14708 11942 14760 11994
rect 14772 11942 14824 11994
rect 14836 11942 14888 11994
rect 23752 11942 23804 11994
rect 23816 11942 23868 11994
rect 23880 11942 23932 11994
rect 23944 11942 23996 11994
rect 2228 11772 2280 11824
rect 3700 11815 3752 11824
rect 3700 11781 3709 11815
rect 3709 11781 3743 11815
rect 3743 11781 3752 11815
rect 3700 11772 3752 11781
rect 4712 11772 4764 11824
rect 6092 11772 6144 11824
rect 6368 11772 6420 11824
rect 8024 11772 8076 11824
rect 10692 11815 10744 11824
rect 10692 11781 10701 11815
rect 10701 11781 10735 11815
rect 10735 11781 10744 11815
rect 10692 11772 10744 11781
rect 12900 11772 12952 11824
rect 9128 11704 9180 11756
rect 13360 11747 13412 11756
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 3148 11679 3200 11688
rect 3148 11645 3157 11679
rect 3157 11645 3191 11679
rect 3191 11645 3200 11679
rect 3148 11636 3200 11645
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 4068 11636 4120 11688
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 3240 11568 3292 11620
rect 6000 11636 6052 11688
rect 8208 11636 8260 11688
rect 8760 11636 8812 11688
rect 10324 11636 10376 11688
rect 5356 11568 5408 11620
rect 7288 11568 7340 11620
rect 4068 11500 4120 11552
rect 5908 11500 5960 11552
rect 12072 11636 12124 11688
rect 12900 11636 12952 11688
rect 11336 11568 11388 11620
rect 11980 11568 12032 11620
rect 12624 11568 12676 11620
rect 13360 11713 13369 11747
rect 13369 11713 13403 11747
rect 13403 11713 13412 11747
rect 13360 11704 13412 11713
rect 13176 11679 13228 11688
rect 13176 11645 13185 11679
rect 13185 11645 13219 11679
rect 13219 11645 13228 11679
rect 13176 11636 13228 11645
rect 13452 11636 13504 11688
rect 14740 11772 14792 11824
rect 14280 11704 14332 11756
rect 15844 11840 15896 11892
rect 21180 11883 21232 11892
rect 16580 11772 16632 11824
rect 16856 11772 16908 11824
rect 13820 11568 13872 11620
rect 14096 11568 14148 11620
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 16948 11636 17000 11688
rect 17132 11636 17184 11688
rect 17960 11636 18012 11688
rect 20260 11704 20312 11756
rect 21180 11849 21189 11883
rect 21189 11849 21223 11883
rect 21223 11849 21232 11883
rect 21180 11840 21232 11849
rect 20720 11772 20772 11824
rect 24584 11840 24636 11892
rect 24860 11883 24912 11892
rect 24860 11849 24869 11883
rect 24869 11849 24903 11883
rect 24903 11849 24912 11883
rect 24860 11840 24912 11849
rect 24952 11840 25004 11892
rect 26148 11840 26200 11892
rect 20076 11679 20128 11688
rect 20076 11645 20085 11679
rect 20085 11645 20119 11679
rect 20119 11645 20128 11679
rect 20076 11636 20128 11645
rect 16580 11568 16632 11620
rect 17408 11568 17460 11620
rect 18052 11568 18104 11620
rect 13084 11500 13136 11552
rect 13544 11500 13596 11552
rect 18144 11500 18196 11552
rect 19616 11500 19668 11552
rect 21548 11704 21600 11756
rect 20628 11679 20680 11688
rect 20628 11645 20637 11679
rect 20637 11645 20671 11679
rect 20671 11645 20680 11679
rect 20628 11636 20680 11645
rect 21180 11636 21232 11688
rect 23480 11636 23532 11688
rect 20812 11611 20864 11620
rect 20812 11577 20821 11611
rect 20821 11577 20855 11611
rect 20855 11577 20864 11611
rect 20812 11568 20864 11577
rect 22100 11568 22152 11620
rect 25504 11636 25556 11688
rect 27252 11704 27304 11756
rect 26516 11636 26568 11688
rect 26240 11611 26292 11620
rect 26240 11577 26249 11611
rect 26249 11577 26283 11611
rect 26283 11577 26292 11611
rect 26240 11568 26292 11577
rect 23296 11543 23348 11552
rect 23296 11509 23305 11543
rect 23305 11509 23339 11543
rect 23339 11509 23348 11543
rect 23296 11500 23348 11509
rect 24400 11500 24452 11552
rect 25596 11500 25648 11552
rect 26608 11543 26660 11552
rect 26608 11509 26617 11543
rect 26617 11509 26651 11543
rect 26651 11509 26660 11543
rect 26608 11500 26660 11509
rect 10090 11398 10142 11450
rect 10154 11398 10206 11450
rect 10218 11398 10270 11450
rect 10282 11398 10334 11450
rect 19198 11398 19250 11450
rect 19262 11398 19314 11450
rect 19326 11398 19378 11450
rect 19390 11398 19442 11450
rect 2136 11296 2188 11348
rect 6000 11296 6052 11348
rect 8208 11296 8260 11348
rect 13544 11296 13596 11348
rect 14280 11296 14332 11348
rect 15384 11296 15436 11348
rect 15568 11296 15620 11348
rect 17408 11296 17460 11348
rect 17960 11296 18012 11348
rect 20628 11296 20680 11348
rect 20996 11296 21048 11348
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 5080 11160 5132 11212
rect 11336 11228 11388 11280
rect 5908 11160 5960 11212
rect 4344 11092 4396 11144
rect 7012 11024 7064 11076
rect 8300 11160 8352 11212
rect 9680 11160 9732 11212
rect 11152 11160 11204 11212
rect 11244 11160 11296 11212
rect 11796 11160 11848 11212
rect 11980 11228 12032 11280
rect 13452 11228 13504 11280
rect 7380 11092 7432 11144
rect 9036 11092 9088 11144
rect 9128 11092 9180 11144
rect 9956 11092 10008 11144
rect 8760 11024 8812 11076
rect 11336 11092 11388 11144
rect 11428 11092 11480 11144
rect 11612 11092 11664 11144
rect 12624 11160 12676 11212
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 15200 11228 15252 11280
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 8484 10956 8536 11008
rect 9496 10956 9548 11008
rect 11244 11024 11296 11076
rect 14372 11092 14424 11144
rect 15384 11160 15436 11212
rect 16488 11228 16540 11280
rect 19892 11228 19944 11280
rect 21456 11228 21508 11280
rect 22192 11228 22244 11280
rect 23480 11296 23532 11348
rect 24584 11296 24636 11348
rect 26332 11296 26384 11348
rect 26516 11296 26568 11348
rect 23112 11228 23164 11280
rect 25596 11271 25648 11280
rect 25596 11237 25605 11271
rect 25605 11237 25639 11271
rect 25639 11237 25648 11271
rect 25596 11228 25648 11237
rect 26608 11271 26660 11280
rect 26608 11237 26642 11271
rect 26642 11237 26660 11271
rect 26608 11228 26660 11237
rect 16764 11203 16816 11212
rect 16764 11169 16773 11203
rect 16773 11169 16807 11203
rect 16807 11169 16816 11203
rect 16764 11160 16816 11169
rect 12164 11024 12216 11076
rect 13176 11024 13228 11076
rect 13636 11024 13688 11076
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 11428 10956 11480 10965
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 12992 10956 13044 11008
rect 15108 11024 15160 11076
rect 15292 10999 15344 11008
rect 15292 10965 15301 10999
rect 15301 10965 15335 10999
rect 15335 10965 15344 10999
rect 15292 10956 15344 10965
rect 16028 11024 16080 11076
rect 16672 11024 16724 11076
rect 16764 11024 16816 11076
rect 17960 11160 18012 11212
rect 18420 11160 18472 11212
rect 20444 11160 20496 11212
rect 20720 11203 20772 11212
rect 17132 11024 17184 11076
rect 19616 11024 19668 11076
rect 19800 11092 19852 11144
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 22652 11203 22704 11212
rect 21548 11024 21600 11076
rect 17408 10956 17460 11008
rect 17592 10956 17644 11008
rect 18420 10956 18472 11008
rect 20904 10956 20956 11008
rect 21916 10956 21968 11008
rect 22652 11169 22661 11203
rect 22661 11169 22695 11203
rect 22695 11169 22704 11203
rect 22652 11160 22704 11169
rect 23756 11203 23808 11212
rect 22744 11024 22796 11076
rect 23020 11024 23072 11076
rect 23756 11169 23765 11203
rect 23765 11169 23799 11203
rect 23799 11169 23808 11203
rect 23756 11160 23808 11169
rect 24124 11203 24176 11212
rect 24124 11169 24133 11203
rect 24133 11169 24167 11203
rect 24167 11169 24176 11203
rect 24124 11160 24176 11169
rect 24952 11160 25004 11212
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 25688 11203 25740 11212
rect 24216 11092 24268 11144
rect 25688 11169 25697 11203
rect 25697 11169 25731 11203
rect 25731 11169 25740 11203
rect 25688 11160 25740 11169
rect 26148 11160 26200 11212
rect 26240 11092 26292 11144
rect 24308 11024 24360 11076
rect 22836 10999 22888 11008
rect 22836 10965 22845 10999
rect 22845 10965 22879 10999
rect 22879 10965 22888 10999
rect 22836 10956 22888 10965
rect 25780 10956 25832 11008
rect 5536 10854 5588 10906
rect 5600 10854 5652 10906
rect 5664 10854 5716 10906
rect 5728 10854 5780 10906
rect 14644 10854 14696 10906
rect 14708 10854 14760 10906
rect 14772 10854 14824 10906
rect 14836 10854 14888 10906
rect 23752 10854 23804 10906
rect 23816 10854 23868 10906
rect 23880 10854 23932 10906
rect 23944 10854 23996 10906
rect 9956 10752 10008 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 4896 10684 4948 10736
rect 1676 10616 1728 10668
rect 4988 10659 5040 10668
rect 2136 10548 2188 10600
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 8208 10684 8260 10736
rect 11336 10684 11388 10736
rect 12348 10752 12400 10804
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 13912 10752 13964 10804
rect 16120 10752 16172 10804
rect 24952 10795 25004 10804
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 3516 10548 3568 10600
rect 4712 10591 4764 10600
rect 4712 10557 4721 10591
rect 4721 10557 4755 10591
rect 4755 10557 4764 10591
rect 4712 10548 4764 10557
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 8024 10616 8076 10668
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 7380 10548 7432 10600
rect 11060 10616 11112 10668
rect 11980 10616 12032 10668
rect 16212 10684 16264 10736
rect 16948 10684 17000 10736
rect 17592 10684 17644 10736
rect 17868 10684 17920 10736
rect 14464 10616 14516 10668
rect 17316 10616 17368 10668
rect 18512 10616 18564 10668
rect 19616 10659 19668 10668
rect 19616 10625 19625 10659
rect 19625 10625 19659 10659
rect 19659 10625 19668 10659
rect 19616 10616 19668 10625
rect 10784 10591 10836 10600
rect 4528 10480 4580 10532
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 9956 10480 10008 10532
rect 11428 10480 11480 10532
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 4252 10412 4304 10464
rect 15292 10548 15344 10600
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 18420 10591 18472 10600
rect 12440 10480 12492 10532
rect 15200 10480 15252 10532
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 18696 10548 18748 10600
rect 20720 10480 20772 10532
rect 25504 10591 25556 10600
rect 23204 10480 23256 10532
rect 25504 10557 25513 10591
rect 25513 10557 25547 10591
rect 25547 10557 25556 10591
rect 25504 10548 25556 10557
rect 25780 10591 25832 10600
rect 25780 10557 25814 10591
rect 25814 10557 25832 10591
rect 25780 10548 25832 10557
rect 26148 10480 26200 10532
rect 12624 10412 12676 10464
rect 13544 10412 13596 10464
rect 15384 10412 15436 10464
rect 16120 10412 16172 10464
rect 18696 10412 18748 10464
rect 20996 10455 21048 10464
rect 20996 10421 21005 10455
rect 21005 10421 21039 10455
rect 21039 10421 21048 10455
rect 20996 10412 21048 10421
rect 22928 10412 22980 10464
rect 24124 10455 24176 10464
rect 24124 10421 24133 10455
rect 24133 10421 24167 10455
rect 24167 10421 24176 10455
rect 24124 10412 24176 10421
rect 25688 10412 25740 10464
rect 10090 10310 10142 10362
rect 10154 10310 10206 10362
rect 10218 10310 10270 10362
rect 10282 10310 10334 10362
rect 19198 10310 19250 10362
rect 19262 10310 19314 10362
rect 19326 10310 19378 10362
rect 19390 10310 19442 10362
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 5908 10208 5960 10260
rect 9956 10208 10008 10260
rect 17684 10208 17736 10260
rect 17868 10208 17920 10260
rect 20444 10208 20496 10260
rect 23480 10208 23532 10260
rect 24216 10251 24268 10260
rect 24216 10217 24225 10251
rect 24225 10217 24259 10251
rect 24259 10217 24268 10251
rect 24216 10208 24268 10217
rect 26148 10208 26200 10260
rect 4804 10140 4856 10192
rect 8300 10140 8352 10192
rect 11980 10140 12032 10192
rect 12532 10140 12584 10192
rect 2688 10072 2740 10124
rect 3516 10072 3568 10124
rect 4988 10072 5040 10124
rect 5908 10072 5960 10124
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 7564 10004 7616 10056
rect 7932 10004 7984 10056
rect 11428 10072 11480 10124
rect 11796 10072 11848 10124
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 17132 10140 17184 10192
rect 12256 10072 12308 10081
rect 17316 10072 17368 10124
rect 11244 10004 11296 10056
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 18880 10072 18932 10124
rect 20536 10072 20588 10124
rect 22836 10140 22888 10192
rect 22928 10140 22980 10192
rect 25504 10140 25556 10192
rect 27528 10183 27580 10192
rect 27528 10149 27537 10183
rect 27537 10149 27571 10183
rect 27571 10149 27580 10183
rect 27528 10140 27580 10149
rect 27804 10140 27856 10192
rect 23572 10072 23624 10124
rect 24124 10115 24176 10124
rect 24124 10081 24133 10115
rect 24133 10081 24167 10115
rect 24167 10081 24176 10115
rect 24124 10072 24176 10081
rect 25596 10115 25648 10124
rect 25596 10081 25630 10115
rect 25630 10081 25648 10115
rect 25596 10072 25648 10081
rect 19892 10004 19944 10056
rect 10324 9936 10376 9988
rect 11612 9936 11664 9988
rect 11704 9936 11756 9988
rect 12256 9936 12308 9988
rect 1676 9868 1728 9920
rect 7564 9868 7616 9920
rect 12532 9868 12584 9920
rect 17592 9868 17644 9920
rect 5536 9766 5588 9818
rect 5600 9766 5652 9818
rect 5664 9766 5716 9818
rect 5728 9766 5780 9818
rect 14644 9766 14696 9818
rect 14708 9766 14760 9818
rect 14772 9766 14824 9818
rect 14836 9766 14888 9818
rect 23752 9766 23804 9818
rect 23816 9766 23868 9818
rect 23880 9766 23932 9818
rect 23944 9766 23996 9818
rect 5908 9707 5960 9716
rect 5908 9673 5917 9707
rect 5917 9673 5951 9707
rect 5951 9673 5960 9707
rect 5908 9664 5960 9673
rect 20628 9664 20680 9716
rect 3148 9596 3200 9648
rect 1676 9528 1728 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 4068 9528 4120 9580
rect 4988 9596 5040 9648
rect 9956 9596 10008 9648
rect 10876 9596 10928 9648
rect 13912 9596 13964 9648
rect 17316 9639 17368 9648
rect 17316 9605 17325 9639
rect 17325 9605 17359 9639
rect 17359 9605 17368 9639
rect 17316 9596 17368 9605
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 5356 9503 5408 9512
rect 2872 9392 2924 9444
rect 2504 9324 2556 9376
rect 4436 9392 4488 9444
rect 3608 9324 3660 9376
rect 4528 9367 4580 9376
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 5540 9435 5592 9444
rect 5540 9401 5549 9435
rect 5549 9401 5583 9435
rect 5583 9401 5592 9435
rect 5540 9392 5592 9401
rect 7564 9460 7616 9512
rect 6736 9392 6788 9444
rect 6920 9392 6972 9444
rect 7472 9392 7524 9444
rect 6644 9324 6696 9376
rect 9404 9460 9456 9512
rect 10692 9460 10744 9512
rect 12164 9460 12216 9512
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 13452 9528 13504 9580
rect 17776 9528 17828 9580
rect 12532 9460 12584 9512
rect 14372 9460 14424 9512
rect 16948 9460 17000 9512
rect 17316 9460 17368 9512
rect 17684 9460 17736 9512
rect 18696 9503 18748 9512
rect 13636 9392 13688 9444
rect 15016 9392 15068 9444
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 19524 9596 19576 9648
rect 19708 9596 19760 9648
rect 20260 9596 20312 9648
rect 20720 9639 20772 9648
rect 20720 9605 20729 9639
rect 20729 9605 20763 9639
rect 20763 9605 20772 9639
rect 20720 9596 20772 9605
rect 19892 9528 19944 9580
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 23296 9571 23348 9580
rect 23296 9537 23305 9571
rect 23305 9537 23339 9571
rect 23339 9537 23348 9571
rect 23296 9528 23348 9537
rect 13728 9324 13780 9376
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 20260 9460 20312 9512
rect 20904 9460 20956 9512
rect 20996 9460 21048 9512
rect 22928 9503 22980 9512
rect 22928 9469 22937 9503
rect 22937 9469 22971 9503
rect 22971 9469 22980 9503
rect 22928 9460 22980 9469
rect 23112 9460 23164 9512
rect 24216 9460 24268 9512
rect 25504 9460 25556 9512
rect 26700 9503 26752 9512
rect 26700 9469 26709 9503
rect 26709 9469 26743 9503
rect 26743 9469 26752 9503
rect 26700 9460 26752 9469
rect 19892 9392 19944 9444
rect 25136 9435 25188 9444
rect 25136 9401 25170 9435
rect 25170 9401 25188 9435
rect 25136 9392 25188 9401
rect 21548 9324 21600 9376
rect 23020 9324 23072 9376
rect 23572 9324 23624 9376
rect 25044 9324 25096 9376
rect 10090 9222 10142 9274
rect 10154 9222 10206 9274
rect 10218 9222 10270 9274
rect 10282 9222 10334 9274
rect 19198 9222 19250 9274
rect 19262 9222 19314 9274
rect 19326 9222 19378 9274
rect 19390 9222 19442 9274
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 4896 9120 4948 9172
rect 5264 9120 5316 9172
rect 6920 9163 6972 9172
rect 2780 9052 2832 9104
rect 3608 9052 3660 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2044 8984 2096 9036
rect 2412 8916 2464 8968
rect 4252 8984 4304 9036
rect 5356 9052 5408 9104
rect 6000 8984 6052 9036
rect 6644 9095 6696 9104
rect 6644 9061 6653 9095
rect 6653 9061 6687 9095
rect 6687 9061 6696 9095
rect 6644 9052 6696 9061
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 7196 9120 7248 9172
rect 7380 9120 7432 9172
rect 7840 9120 7892 9172
rect 7472 9052 7524 9104
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 7196 8984 7248 9036
rect 9128 9052 9180 9104
rect 9220 8984 9272 9036
rect 9634 9052 9686 9104
rect 10416 9120 10468 9172
rect 10784 9120 10836 9172
rect 13728 9120 13780 9172
rect 20536 9163 20588 9172
rect 20536 9129 20545 9163
rect 20545 9129 20579 9163
rect 20579 9129 20588 9163
rect 20536 9120 20588 9129
rect 23204 9120 23256 9172
rect 24216 9163 24268 9172
rect 24216 9129 24225 9163
rect 24225 9129 24259 9163
rect 24259 9129 24268 9163
rect 24216 9120 24268 9129
rect 25596 9120 25648 9172
rect 26424 9120 26476 9172
rect 7840 8916 7892 8968
rect 10048 8984 10100 9036
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 11060 9027 11112 9036
rect 11060 8993 11069 9027
rect 11069 8993 11103 9027
rect 11103 8993 11112 9027
rect 11060 8984 11112 8993
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 11612 8984 11664 9036
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 15016 9095 15068 9104
rect 12900 8984 12952 9036
rect 13452 8984 13504 9036
rect 10416 8916 10468 8968
rect 13636 8916 13688 8968
rect 4988 8848 5040 8900
rect 5356 8848 5408 8900
rect 15016 9061 15025 9095
rect 15025 9061 15059 9095
rect 15059 9061 15068 9095
rect 15016 9052 15068 9061
rect 15660 9052 15712 9104
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 16304 8984 16356 9036
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 16948 8984 17000 9036
rect 17224 9052 17276 9104
rect 17776 9052 17828 9104
rect 19892 9052 19944 9104
rect 20444 9052 20496 9104
rect 22100 9052 22152 9104
rect 19800 8984 19852 9036
rect 15752 8916 15804 8968
rect 19892 8916 19944 8968
rect 17592 8848 17644 8900
rect 17868 8891 17920 8900
rect 17868 8857 17877 8891
rect 17877 8857 17911 8891
rect 17911 8857 17920 8891
rect 17868 8848 17920 8857
rect 5908 8780 5960 8832
rect 8484 8780 8536 8832
rect 10784 8780 10836 8832
rect 11612 8780 11664 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 12900 8780 12952 8832
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 16856 8780 16908 8832
rect 17776 8780 17828 8832
rect 19708 8848 19760 8900
rect 21824 8984 21876 9036
rect 23020 9027 23072 9036
rect 23020 8993 23029 9027
rect 23029 8993 23063 9027
rect 23063 8993 23072 9027
rect 23020 8984 23072 8993
rect 21916 8916 21968 8968
rect 25044 8984 25096 9036
rect 25320 8984 25372 9036
rect 26148 9052 26200 9104
rect 26792 9027 26844 9036
rect 25412 8916 25464 8968
rect 21824 8848 21876 8900
rect 26792 8993 26801 9027
rect 26801 8993 26835 9027
rect 26835 8993 26844 9027
rect 26792 8984 26844 8993
rect 27528 9027 27580 9036
rect 27528 8993 27537 9027
rect 27537 8993 27571 9027
rect 27571 8993 27580 9027
rect 27528 8984 27580 8993
rect 27712 8891 27764 8900
rect 27712 8857 27721 8891
rect 27721 8857 27755 8891
rect 27755 8857 27764 8891
rect 27712 8848 27764 8857
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 18696 8780 18748 8832
rect 19616 8780 19668 8832
rect 22008 8780 22060 8832
rect 24952 8780 25004 8832
rect 5536 8678 5588 8730
rect 5600 8678 5652 8730
rect 5664 8678 5716 8730
rect 5728 8678 5780 8730
rect 14644 8678 14696 8730
rect 14708 8678 14760 8730
rect 14772 8678 14824 8730
rect 14836 8678 14888 8730
rect 23752 8678 23804 8730
rect 23816 8678 23868 8730
rect 23880 8678 23932 8730
rect 23944 8678 23996 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 4160 8576 4212 8628
rect 4712 8576 4764 8628
rect 7840 8576 7892 8628
rect 5172 8508 5224 8560
rect 10048 8576 10100 8628
rect 9220 8508 9272 8560
rect 11336 8576 11388 8628
rect 15752 8619 15804 8628
rect 2412 8440 2464 8492
rect 2044 8372 2096 8424
rect 2504 8415 2556 8424
rect 2504 8381 2513 8415
rect 2513 8381 2547 8415
rect 2547 8381 2556 8415
rect 2504 8372 2556 8381
rect 9404 8440 9456 8492
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8300 8372 8352 8424
rect 8484 8415 8536 8424
rect 8484 8381 8518 8415
rect 8518 8381 8536 8415
rect 8484 8372 8536 8381
rect 9680 8372 9732 8424
rect 10784 8372 10836 8424
rect 12072 8415 12124 8424
rect 3608 8304 3660 8356
rect 8760 8304 8812 8356
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 12164 8372 12216 8424
rect 12532 8372 12584 8424
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 18972 8576 19024 8628
rect 20168 8619 20220 8628
rect 20168 8585 20177 8619
rect 20177 8585 20211 8619
rect 20211 8585 20220 8619
rect 20168 8576 20220 8585
rect 22744 8576 22796 8628
rect 23204 8576 23256 8628
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 17776 8508 17828 8560
rect 20260 8508 20312 8560
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 20076 8440 20128 8492
rect 15568 8372 15620 8424
rect 17224 8372 17276 8424
rect 18052 8372 18104 8424
rect 18696 8372 18748 8424
rect 19064 8415 19116 8424
rect 19064 8381 19098 8415
rect 19098 8381 19116 8415
rect 19064 8372 19116 8381
rect 20168 8372 20220 8424
rect 21732 8372 21784 8424
rect 23480 8372 23532 8424
rect 24400 8372 24452 8424
rect 25320 8508 25372 8560
rect 26240 8508 26292 8560
rect 25044 8440 25096 8492
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 25136 8372 25188 8424
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 26700 8415 26752 8424
rect 11060 8304 11112 8356
rect 11980 8304 12032 8356
rect 13544 8347 13596 8356
rect 13544 8313 13553 8347
rect 13553 8313 13587 8347
rect 13587 8313 13596 8347
rect 13544 8304 13596 8313
rect 14188 8304 14240 8356
rect 17592 8304 17644 8356
rect 7012 8236 7064 8288
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 18696 8236 18748 8288
rect 20720 8236 20772 8288
rect 21180 8236 21232 8288
rect 22192 8304 22244 8356
rect 23112 8236 23164 8288
rect 24952 8236 25004 8288
rect 25504 8236 25556 8288
rect 25596 8236 25648 8288
rect 26700 8381 26709 8415
rect 26709 8381 26743 8415
rect 26743 8381 26752 8415
rect 26700 8372 26752 8381
rect 26884 8279 26936 8288
rect 26884 8245 26893 8279
rect 26893 8245 26927 8279
rect 26927 8245 26936 8279
rect 26884 8236 26936 8245
rect 10090 8134 10142 8186
rect 10154 8134 10206 8186
rect 10218 8134 10270 8186
rect 10282 8134 10334 8186
rect 19198 8134 19250 8186
rect 19262 8134 19314 8186
rect 19326 8134 19378 8186
rect 19390 8134 19442 8186
rect 1492 8032 1544 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 1584 7896 1636 7948
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 5080 7896 5132 7948
rect 5172 7828 5224 7880
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 8300 8032 8352 8084
rect 12164 8032 12216 8084
rect 15476 8032 15528 8084
rect 12624 8007 12676 8016
rect 5448 7896 5500 7905
rect 6000 7896 6052 7948
rect 6092 7896 6144 7948
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 7840 7828 7892 7880
rect 9956 7896 10008 7948
rect 11336 7896 11388 7948
rect 12624 7973 12658 8007
rect 12658 7973 12676 8007
rect 12624 7964 12676 7973
rect 15292 7964 15344 8016
rect 18512 8032 18564 8084
rect 18972 8032 19024 8084
rect 21088 8032 21140 8084
rect 22928 8032 22980 8084
rect 13084 7896 13136 7948
rect 14372 7896 14424 7948
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 17684 7939 17736 7948
rect 17684 7905 17693 7939
rect 17693 7905 17727 7939
rect 17727 7905 17736 7939
rect 17684 7896 17736 7905
rect 17132 7828 17184 7880
rect 17868 7939 17920 7948
rect 17868 7905 17877 7939
rect 17877 7905 17911 7939
rect 17911 7905 17920 7939
rect 18512 7939 18564 7948
rect 17868 7896 17920 7905
rect 18512 7905 18521 7939
rect 18521 7905 18555 7939
rect 18555 7905 18564 7939
rect 18512 7896 18564 7905
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 18052 7828 18104 7880
rect 18972 7896 19024 7948
rect 20076 7896 20128 7948
rect 21824 7964 21876 8016
rect 25780 8032 25832 8084
rect 25964 8032 26016 8084
rect 26240 8007 26292 8016
rect 20904 7896 20956 7948
rect 21180 7896 21232 7948
rect 22100 7896 22152 7948
rect 22836 7939 22888 7948
rect 20168 7828 20220 7880
rect 16396 7760 16448 7812
rect 21272 7828 21324 7880
rect 22836 7905 22845 7939
rect 22845 7905 22879 7939
rect 22879 7905 22888 7939
rect 22836 7896 22888 7905
rect 23020 7939 23072 7948
rect 23020 7905 23029 7939
rect 23029 7905 23063 7939
rect 23063 7905 23072 7939
rect 23020 7896 23072 7905
rect 26240 7973 26274 8007
rect 26274 7973 26292 8007
rect 26240 7964 26292 7973
rect 22744 7828 22796 7880
rect 24860 7896 24912 7948
rect 25504 7896 25556 7948
rect 24952 7828 25004 7880
rect 11152 7692 11204 7744
rect 12256 7692 12308 7744
rect 16304 7692 16356 7744
rect 17776 7692 17828 7744
rect 17960 7692 18012 7744
rect 19064 7735 19116 7744
rect 19064 7701 19073 7735
rect 19073 7701 19107 7735
rect 19107 7701 19116 7735
rect 19064 7692 19116 7701
rect 22836 7692 22888 7744
rect 24216 7692 24268 7744
rect 24768 7692 24820 7744
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 5536 7590 5588 7642
rect 5600 7590 5652 7642
rect 5664 7590 5716 7642
rect 5728 7590 5780 7642
rect 14644 7590 14696 7642
rect 14708 7590 14760 7642
rect 14772 7590 14824 7642
rect 14836 7590 14888 7642
rect 23752 7590 23804 7642
rect 23816 7590 23868 7642
rect 23880 7590 23932 7642
rect 23944 7590 23996 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 4068 7488 4120 7540
rect 3976 7463 4028 7472
rect 3976 7429 3985 7463
rect 3985 7429 4019 7463
rect 4019 7429 4028 7463
rect 3976 7420 4028 7429
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 2412 7352 2464 7404
rect 4160 7352 4212 7404
rect 5356 7488 5408 7540
rect 6000 7488 6052 7540
rect 6828 7488 6880 7540
rect 10876 7488 10928 7540
rect 11888 7488 11940 7540
rect 17040 7488 17092 7540
rect 17316 7488 17368 7540
rect 19708 7531 19760 7540
rect 8116 7420 8168 7472
rect 12808 7420 12860 7472
rect 13268 7420 13320 7472
rect 5908 7352 5960 7404
rect 7196 7352 7248 7404
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 2872 7284 2924 7336
rect 3148 7216 3200 7268
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 4068 7284 4120 7336
rect 4988 7284 5040 7336
rect 5172 7284 5224 7336
rect 6552 7284 6604 7336
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 7656 7352 7708 7404
rect 8392 7352 8444 7404
rect 7840 7327 7892 7336
rect 5908 7216 5960 7268
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 13360 7352 13412 7404
rect 17592 7352 17644 7404
rect 19708 7497 19717 7531
rect 19717 7497 19751 7531
rect 19751 7497 19760 7531
rect 19708 7488 19760 7497
rect 20076 7531 20128 7540
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 23388 7488 23440 7540
rect 23480 7488 23532 7540
rect 18972 7420 19024 7472
rect 21180 7352 21232 7404
rect 12164 7284 12216 7336
rect 12256 7284 12308 7336
rect 16488 7284 16540 7336
rect 17960 7327 18012 7336
rect 17960 7293 17994 7327
rect 17994 7293 18012 7327
rect 17960 7284 18012 7293
rect 19984 7284 20036 7336
rect 20536 7284 20588 7336
rect 21824 7352 21876 7404
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 23020 7352 23072 7404
rect 23480 7352 23532 7404
rect 21456 7327 21508 7336
rect 21456 7293 21465 7327
rect 21465 7293 21499 7327
rect 21499 7293 21508 7327
rect 21456 7284 21508 7293
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 22652 7284 22704 7336
rect 23112 7327 23164 7336
rect 23112 7293 23121 7327
rect 23121 7293 23155 7327
rect 23155 7293 23164 7327
rect 23112 7284 23164 7293
rect 22100 7216 22152 7268
rect 22836 7216 22888 7268
rect 4712 7148 4764 7200
rect 7380 7148 7432 7200
rect 8024 7148 8076 7200
rect 18052 7148 18104 7200
rect 22468 7148 22520 7200
rect 23848 7327 23900 7336
rect 23848 7293 23857 7327
rect 23857 7293 23891 7327
rect 23891 7293 23900 7327
rect 23848 7284 23900 7293
rect 24860 7327 24912 7336
rect 24032 7259 24084 7268
rect 24032 7225 24041 7259
rect 24041 7225 24075 7259
rect 24075 7225 24084 7259
rect 24032 7216 24084 7225
rect 24860 7293 24869 7327
rect 24869 7293 24903 7327
rect 24903 7293 24912 7327
rect 24860 7284 24912 7293
rect 25596 7284 25648 7336
rect 10090 7046 10142 7098
rect 10154 7046 10206 7098
rect 10218 7046 10270 7098
rect 10282 7046 10334 7098
rect 19198 7046 19250 7098
rect 19262 7046 19314 7098
rect 19326 7046 19378 7098
rect 19390 7046 19442 7098
rect 4068 6944 4120 6996
rect 2688 6876 2740 6928
rect 2412 6808 2464 6860
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 4712 6808 4764 6860
rect 6184 6851 6236 6860
rect 5356 6740 5408 6792
rect 4252 6672 4304 6724
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 6644 6808 6696 6860
rect 7380 6851 7432 6860
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 7656 6876 7708 6928
rect 11336 6944 11388 6996
rect 18512 6944 18564 6996
rect 23848 6944 23900 6996
rect 24860 6944 24912 6996
rect 26056 6944 26108 6996
rect 11152 6919 11204 6928
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 11152 6885 11161 6919
rect 11161 6885 11195 6919
rect 11195 6885 11204 6919
rect 11152 6876 11204 6885
rect 10876 6851 10928 6860
rect 9680 6740 9732 6792
rect 7288 6672 7340 6724
rect 8116 6672 8168 6724
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 10508 6740 10560 6792
rect 10692 6740 10744 6792
rect 12440 6808 12492 6860
rect 17592 6876 17644 6928
rect 20260 6919 20312 6928
rect 16396 6808 16448 6860
rect 16948 6808 17000 6860
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 20260 6885 20269 6919
rect 20269 6885 20303 6919
rect 20303 6885 20312 6919
rect 20260 6876 20312 6885
rect 18788 6808 18840 6860
rect 21088 6851 21140 6860
rect 21088 6817 21122 6851
rect 21122 6817 21140 6851
rect 22468 6876 22520 6928
rect 25136 6876 25188 6928
rect 25504 6919 25556 6928
rect 11796 6740 11848 6792
rect 21088 6808 21140 6817
rect 23204 6808 23256 6860
rect 24584 6808 24636 6860
rect 25504 6885 25513 6919
rect 25513 6885 25547 6919
rect 25547 6885 25556 6919
rect 25504 6876 25556 6885
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 25596 6851 25648 6860
rect 25596 6817 25605 6851
rect 25605 6817 25639 6851
rect 25639 6817 25648 6851
rect 25596 6808 25648 6817
rect 11888 6672 11940 6724
rect 17868 6672 17920 6724
rect 22468 6740 22520 6792
rect 23664 6672 23716 6724
rect 26056 6740 26108 6792
rect 2136 6604 2188 6656
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 3424 6604 3476 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7012 6604 7064 6656
rect 7472 6604 7524 6656
rect 10140 6604 10192 6656
rect 12992 6604 13044 6656
rect 16488 6604 16540 6656
rect 20812 6604 20864 6656
rect 22836 6604 22888 6656
rect 26884 6604 26936 6656
rect 5536 6502 5588 6554
rect 5600 6502 5652 6554
rect 5664 6502 5716 6554
rect 5728 6502 5780 6554
rect 14644 6502 14696 6554
rect 14708 6502 14760 6554
rect 14772 6502 14824 6554
rect 14836 6502 14888 6554
rect 23752 6502 23804 6554
rect 23816 6502 23868 6554
rect 23880 6502 23932 6554
rect 23944 6502 23996 6554
rect 3240 6400 3292 6452
rect 4068 6400 4120 6452
rect 6644 6400 6696 6452
rect 8116 6400 8168 6452
rect 10784 6400 10836 6452
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 17684 6443 17736 6452
rect 17684 6409 17693 6443
rect 17693 6409 17727 6443
rect 17727 6409 17736 6443
rect 17684 6400 17736 6409
rect 21088 6443 21140 6452
rect 21088 6409 21097 6443
rect 21097 6409 21131 6443
rect 21131 6409 21140 6443
rect 21088 6400 21140 6409
rect 5356 6332 5408 6384
rect 23572 6400 23624 6452
rect 24308 6400 24360 6452
rect 22836 6332 22888 6384
rect 24584 6400 24636 6452
rect 4252 6264 4304 6316
rect 12256 6264 12308 6316
rect 17316 6264 17368 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2136 6128 2188 6180
rect 3424 6196 3476 6248
rect 7012 6196 7064 6248
rect 7656 6196 7708 6248
rect 8484 6239 8536 6248
rect 4068 6128 4120 6180
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 8392 6128 8444 6180
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 10508 6196 10560 6248
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 14004 6239 14056 6248
rect 9496 6060 9548 6112
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 15200 6196 15252 6248
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 16396 6196 16448 6248
rect 17408 6196 17460 6248
rect 17868 6196 17920 6248
rect 20536 6239 20588 6248
rect 13728 6128 13780 6180
rect 14648 6128 14700 6180
rect 16488 6128 16540 6180
rect 16948 6128 17000 6180
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 22928 6264 22980 6316
rect 21272 6196 21324 6248
rect 23112 6239 23164 6248
rect 23112 6205 23121 6239
rect 23121 6205 23155 6239
rect 23155 6205 23164 6239
rect 23112 6196 23164 6205
rect 23572 6196 23624 6248
rect 24308 6239 24360 6248
rect 24308 6205 24317 6239
rect 24317 6205 24351 6239
rect 24351 6205 24360 6239
rect 24308 6196 24360 6205
rect 26148 6196 26200 6248
rect 25320 6128 25372 6180
rect 14464 6060 14516 6112
rect 15016 6060 15068 6112
rect 15936 6060 15988 6112
rect 16856 6060 16908 6112
rect 22100 6060 22152 6112
rect 23296 6060 23348 6112
rect 23664 6060 23716 6112
rect 24676 6060 24728 6112
rect 24768 6103 24820 6112
rect 24768 6069 24777 6103
rect 24777 6069 24811 6103
rect 24811 6069 24820 6103
rect 24768 6060 24820 6069
rect 10090 5958 10142 6010
rect 10154 5958 10206 6010
rect 10218 5958 10270 6010
rect 10282 5958 10334 6010
rect 19198 5958 19250 6010
rect 19262 5958 19314 6010
rect 19326 5958 19378 6010
rect 19390 5958 19442 6010
rect 5908 5856 5960 5908
rect 7840 5856 7892 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 9864 5856 9916 5908
rect 10508 5856 10560 5908
rect 12624 5856 12676 5908
rect 12900 5856 12952 5908
rect 16580 5856 16632 5908
rect 3148 5720 3200 5772
rect 8300 5720 8352 5772
rect 10416 5788 10468 5840
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 9588 5652 9640 5704
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 10508 5763 10560 5772
rect 9864 5720 9916 5729
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 10876 5720 10928 5772
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 9956 5652 10008 5704
rect 11796 5720 11848 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 13820 5788 13872 5840
rect 14004 5720 14056 5772
rect 15108 5788 15160 5840
rect 17408 5788 17460 5840
rect 20536 5788 20588 5840
rect 22560 5856 22612 5908
rect 22744 5856 22796 5908
rect 23388 5856 23440 5908
rect 24860 5856 24912 5908
rect 16212 5720 16264 5772
rect 16948 5720 17000 5772
rect 19800 5720 19852 5772
rect 20444 5720 20496 5772
rect 12440 5652 12492 5704
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 15292 5652 15344 5704
rect 16488 5652 16540 5704
rect 18420 5652 18472 5704
rect 1860 5516 1912 5568
rect 14648 5584 14700 5636
rect 24400 5788 24452 5840
rect 27436 5788 27488 5840
rect 27712 5831 27764 5840
rect 27712 5797 27721 5831
rect 27721 5797 27755 5831
rect 27755 5797 27764 5831
rect 27712 5788 27764 5797
rect 22744 5720 22796 5772
rect 23664 5763 23716 5772
rect 23664 5729 23673 5763
rect 23673 5729 23707 5763
rect 23707 5729 23716 5763
rect 23664 5720 23716 5729
rect 23020 5652 23072 5704
rect 9680 5516 9732 5568
rect 10876 5516 10928 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 17224 5516 17276 5568
rect 19616 5516 19668 5568
rect 27160 5584 27212 5636
rect 22836 5559 22888 5568
rect 22836 5525 22845 5559
rect 22845 5525 22879 5559
rect 22879 5525 22888 5559
rect 22836 5516 22888 5525
rect 24124 5516 24176 5568
rect 5536 5414 5588 5466
rect 5600 5414 5652 5466
rect 5664 5414 5716 5466
rect 5728 5414 5780 5466
rect 14644 5414 14696 5466
rect 14708 5414 14760 5466
rect 14772 5414 14824 5466
rect 14836 5414 14888 5466
rect 23752 5414 23804 5466
rect 23816 5414 23868 5466
rect 23880 5414 23932 5466
rect 23944 5414 23996 5466
rect 3884 5312 3936 5364
rect 7748 5312 7800 5364
rect 7656 5244 7708 5296
rect 9496 5244 9548 5296
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 8300 5176 8352 5228
rect 9772 5176 9824 5228
rect 22284 5312 22336 5364
rect 22468 5312 22520 5364
rect 22836 5312 22888 5364
rect 23388 5312 23440 5364
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 12532 5244 12584 5296
rect 14464 5244 14516 5296
rect 16212 5244 16264 5296
rect 17684 5244 17736 5296
rect 21548 5287 21600 5296
rect 14096 5176 14148 5228
rect 12072 5151 12124 5160
rect 2780 5040 2832 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 9956 5040 10008 5092
rect 9864 4972 9916 5024
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 12532 5108 12584 5160
rect 12808 5108 12860 5160
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 10508 5083 10560 5092
rect 10508 5049 10517 5083
rect 10517 5049 10551 5083
rect 10551 5049 10560 5083
rect 10508 5040 10560 5049
rect 11428 5040 11480 5092
rect 12256 5083 12308 5092
rect 12256 5049 12265 5083
rect 12265 5049 12299 5083
rect 12299 5049 12308 5083
rect 12256 5040 12308 5049
rect 12072 4972 12124 5024
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 13452 5040 13504 5092
rect 13544 4972 13596 5024
rect 17960 5176 18012 5228
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16488 5108 16540 5160
rect 17408 5151 17460 5160
rect 17408 5117 17417 5151
rect 17417 5117 17451 5151
rect 17451 5117 17460 5151
rect 17408 5108 17460 5117
rect 18144 5176 18196 5228
rect 21548 5253 21557 5287
rect 21557 5253 21591 5287
rect 21591 5253 21600 5287
rect 21548 5244 21600 5253
rect 24400 5312 24452 5364
rect 18420 5151 18472 5160
rect 18420 5117 18429 5151
rect 18429 5117 18463 5151
rect 18463 5117 18472 5151
rect 18420 5108 18472 5117
rect 18696 5108 18748 5160
rect 20996 5108 21048 5160
rect 16580 5040 16632 5092
rect 18236 5083 18288 5092
rect 18236 5049 18245 5083
rect 18245 5049 18279 5083
rect 18279 5049 18288 5083
rect 18236 5040 18288 5049
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 15108 4972 15160 5024
rect 19064 4972 19116 5024
rect 19524 5040 19576 5092
rect 22100 5040 22152 5092
rect 22744 5108 22796 5160
rect 22928 5151 22980 5160
rect 22928 5117 22937 5151
rect 22937 5117 22971 5151
rect 22971 5117 22980 5151
rect 22928 5108 22980 5117
rect 23020 5151 23072 5160
rect 23020 5117 23029 5151
rect 23029 5117 23063 5151
rect 23063 5117 23072 5151
rect 27620 5176 27672 5228
rect 23020 5108 23072 5117
rect 22376 5040 22428 5092
rect 26884 5108 26936 5160
rect 19984 4972 20036 5024
rect 20444 5015 20496 5024
rect 20444 4981 20453 5015
rect 20453 4981 20487 5015
rect 20487 4981 20496 5015
rect 20444 4972 20496 4981
rect 22284 4972 22336 5024
rect 24124 5040 24176 5092
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 24400 4972 24452 5024
rect 10090 4870 10142 4922
rect 10154 4870 10206 4922
rect 10218 4870 10270 4922
rect 10282 4870 10334 4922
rect 19198 4870 19250 4922
rect 19262 4870 19314 4922
rect 19326 4870 19378 4922
rect 19390 4870 19442 4922
rect 1584 4768 1636 4820
rect 1768 4700 1820 4752
rect 2412 4700 2464 4752
rect 3884 4700 3936 4752
rect 2504 4675 2556 4684
rect 2504 4641 2513 4675
rect 2513 4641 2547 4675
rect 2547 4641 2556 4675
rect 2504 4632 2556 4641
rect 2872 4632 2924 4684
rect 4896 4632 4948 4684
rect 4160 4564 4212 4616
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 6920 4768 6972 4820
rect 9128 4768 9180 4820
rect 9956 4768 10008 4820
rect 10692 4768 10744 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 6184 4632 6236 4684
rect 8484 4632 8536 4684
rect 9680 4700 9732 4752
rect 9772 4743 9824 4752
rect 9772 4709 9781 4743
rect 9781 4709 9815 4743
rect 9815 4709 9824 4743
rect 9772 4700 9824 4709
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 11796 4700 11848 4752
rect 12256 4700 12308 4752
rect 15016 4743 15068 4752
rect 15016 4709 15050 4743
rect 15050 4709 15068 4743
rect 15016 4700 15068 4709
rect 16948 4700 17000 4752
rect 19708 4700 19760 4752
rect 20260 4743 20312 4752
rect 20260 4709 20269 4743
rect 20269 4709 20303 4743
rect 20303 4709 20312 4743
rect 20628 4768 20680 4820
rect 20996 4811 21048 4820
rect 20996 4777 21005 4811
rect 21005 4777 21039 4811
rect 21039 4777 21048 4811
rect 20996 4768 21048 4777
rect 22928 4768 22980 4820
rect 20260 4700 20312 4709
rect 12808 4632 12860 4684
rect 2780 4496 2832 4548
rect 2964 4428 3016 4480
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 12164 4564 12216 4616
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 15292 4632 15344 4684
rect 17684 4675 17736 4684
rect 17684 4641 17693 4675
rect 17693 4641 17727 4675
rect 17727 4641 17736 4675
rect 17684 4632 17736 4641
rect 17776 4632 17828 4684
rect 20168 4675 20220 4684
rect 20168 4641 20177 4675
rect 20177 4641 20211 4675
rect 20211 4641 20220 4675
rect 20168 4632 20220 4641
rect 21180 4675 21232 4684
rect 18696 4564 18748 4616
rect 21180 4641 21189 4675
rect 21189 4641 21223 4675
rect 21223 4641 21232 4675
rect 21180 4632 21232 4641
rect 23204 4700 23256 4752
rect 27528 4743 27580 4752
rect 27528 4709 27537 4743
rect 27537 4709 27571 4743
rect 27571 4709 27580 4743
rect 27528 4700 27580 4709
rect 25412 4675 25464 4684
rect 14464 4496 14516 4548
rect 17224 4539 17276 4548
rect 17224 4505 17233 4539
rect 17233 4505 17267 4539
rect 17267 4505 17276 4539
rect 17224 4496 17276 4505
rect 18972 4496 19024 4548
rect 14096 4428 14148 4480
rect 14372 4428 14424 4480
rect 18052 4428 18104 4480
rect 20260 4428 20312 4480
rect 20352 4428 20404 4480
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 25412 4641 25421 4675
rect 25421 4641 25455 4675
rect 25455 4641 25464 4675
rect 25412 4632 25464 4641
rect 26056 4632 26108 4684
rect 26792 4675 26844 4684
rect 26792 4641 26801 4675
rect 26801 4641 26835 4675
rect 26835 4641 26844 4675
rect 26792 4632 26844 4641
rect 24216 4496 24268 4548
rect 25228 4471 25280 4480
rect 25228 4437 25237 4471
rect 25237 4437 25271 4471
rect 25271 4437 25280 4471
rect 25228 4428 25280 4437
rect 26332 4471 26384 4480
rect 26332 4437 26341 4471
rect 26341 4437 26375 4471
rect 26375 4437 26384 4471
rect 26332 4428 26384 4437
rect 5536 4326 5588 4378
rect 5600 4326 5652 4378
rect 5664 4326 5716 4378
rect 5728 4326 5780 4378
rect 14644 4326 14696 4378
rect 14708 4326 14760 4378
rect 14772 4326 14824 4378
rect 14836 4326 14888 4378
rect 23752 4326 23804 4378
rect 23816 4326 23868 4378
rect 23880 4326 23932 4378
rect 23944 4326 23996 4378
rect 2504 4267 2556 4276
rect 2504 4233 2513 4267
rect 2513 4233 2547 4267
rect 2547 4233 2556 4267
rect 2504 4224 2556 4233
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 10508 4224 10560 4276
rect 2780 4020 2832 4072
rect 3148 4063 3200 4072
rect 3148 4029 3157 4063
rect 3157 4029 3191 4063
rect 3191 4029 3200 4063
rect 3148 4020 3200 4029
rect 4252 4020 4304 4072
rect 6184 4088 6236 4140
rect 8300 4088 8352 4140
rect 10416 4088 10468 4140
rect 12440 4224 12492 4276
rect 12808 4224 12860 4276
rect 13544 4224 13596 4276
rect 13360 4156 13412 4208
rect 18236 4224 18288 4276
rect 26332 4224 26384 4276
rect 13084 4088 13136 4140
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 15292 4156 15344 4208
rect 17684 4156 17736 4208
rect 18144 4088 18196 4140
rect 18328 4156 18380 4208
rect 18972 4156 19024 4208
rect 19984 4156 20036 4208
rect 18420 4088 18472 4140
rect 2872 3952 2924 4004
rect 1400 3884 1452 3936
rect 2596 3884 2648 3936
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 5356 4063 5408 4072
rect 4712 4020 4764 4029
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 4528 3995 4580 4004
rect 4528 3961 4537 3995
rect 4537 3961 4571 3995
rect 4571 3961 4580 3995
rect 4528 3952 4580 3961
rect 9496 4020 9548 4072
rect 12164 4020 12216 4072
rect 12624 4020 12676 4072
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14096 4020 14148 4072
rect 5356 3884 5408 3936
rect 7104 3952 7156 4004
rect 7196 3952 7248 4004
rect 9680 3952 9732 4004
rect 9864 3952 9916 4004
rect 12532 3952 12584 4004
rect 13360 3952 13412 4004
rect 16948 4020 17000 4072
rect 17960 4063 18012 4072
rect 17960 4029 17969 4063
rect 17969 4029 18003 4063
rect 18003 4029 18012 4063
rect 17960 4020 18012 4029
rect 18696 4020 18748 4072
rect 20720 4088 20772 4140
rect 21640 4088 21692 4140
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 19064 4020 19116 4072
rect 21088 4020 21140 4072
rect 22008 4020 22060 4072
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 23388 4020 23440 4072
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 25964 4063 26016 4072
rect 25964 4029 25973 4063
rect 25973 4029 26007 4063
rect 26007 4029 26016 4063
rect 25964 4020 26016 4029
rect 15108 3952 15160 4004
rect 16672 3952 16724 4004
rect 5724 3884 5776 3936
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 7932 3884 7984 3936
rect 12992 3884 13044 3936
rect 13176 3884 13228 3936
rect 14096 3884 14148 3936
rect 16120 3884 16172 3936
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 18328 3884 18380 3936
rect 19524 3884 19576 3936
rect 20168 3884 20220 3936
rect 22652 3884 22704 3936
rect 23388 3884 23440 3936
rect 23940 3952 23992 4004
rect 27620 3952 27672 4004
rect 24952 3884 25004 3936
rect 26148 3927 26200 3936
rect 26148 3893 26157 3927
rect 26157 3893 26191 3927
rect 26191 3893 26200 3927
rect 26148 3884 26200 3893
rect 10090 3782 10142 3834
rect 10154 3782 10206 3834
rect 10218 3782 10270 3834
rect 10282 3782 10334 3834
rect 19198 3782 19250 3834
rect 19262 3782 19314 3834
rect 19326 3782 19378 3834
rect 19390 3782 19442 3834
rect 5724 3680 5776 3732
rect 5908 3612 5960 3664
rect 7104 3680 7156 3732
rect 9588 3612 9640 3664
rect 1492 3587 1544 3596
rect 1492 3553 1501 3587
rect 1501 3553 1535 3587
rect 1535 3553 1544 3587
rect 1492 3544 1544 3553
rect 1768 3544 1820 3596
rect 2320 3544 2372 3596
rect 4804 3544 4856 3596
rect 7840 3544 7892 3596
rect 8760 3544 8812 3596
rect 9864 3544 9916 3596
rect 8668 3476 8720 3528
rect 9680 3476 9732 3528
rect 9772 3476 9824 3528
rect 10692 3544 10744 3596
rect 12440 3612 12492 3664
rect 12900 3680 12952 3732
rect 19708 3680 19760 3732
rect 21180 3680 21232 3732
rect 23020 3680 23072 3732
rect 23848 3680 23900 3732
rect 12716 3544 12768 3596
rect 11980 3476 12032 3528
rect 13912 3612 13964 3664
rect 14372 3612 14424 3664
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 13268 3544 13320 3596
rect 15660 3544 15712 3596
rect 16764 3544 16816 3596
rect 15292 3476 15344 3528
rect 18236 3612 18288 3664
rect 20444 3612 20496 3664
rect 22008 3612 22060 3664
rect 22744 3612 22796 3664
rect 17040 3544 17092 3596
rect 18052 3544 18104 3596
rect 18880 3587 18932 3596
rect 18880 3553 18889 3587
rect 18889 3553 18923 3587
rect 18923 3553 18932 3587
rect 18880 3544 18932 3553
rect 19984 3587 20036 3596
rect 19984 3553 19993 3587
rect 19993 3553 20027 3587
rect 20027 3553 20036 3587
rect 19984 3544 20036 3553
rect 20536 3544 20588 3596
rect 20260 3476 20312 3528
rect 21272 3544 21324 3596
rect 23388 3544 23440 3596
rect 25228 3612 25280 3664
rect 25688 3612 25740 3664
rect 26516 3612 26568 3664
rect 9496 3408 9548 3460
rect 940 3340 992 3392
rect 4068 3340 4120 3392
rect 6552 3340 6604 3392
rect 8668 3340 8720 3392
rect 10508 3383 10560 3392
rect 10508 3349 10517 3383
rect 10517 3349 10551 3383
rect 10551 3349 10560 3383
rect 10508 3340 10560 3349
rect 12532 3408 12584 3460
rect 13176 3408 13228 3460
rect 15476 3408 15528 3460
rect 23848 3587 23900 3596
rect 23848 3553 23857 3587
rect 23857 3553 23891 3587
rect 23891 3553 23900 3587
rect 23848 3544 23900 3553
rect 24400 3544 24452 3596
rect 25412 3544 25464 3596
rect 26424 3544 26476 3596
rect 27068 3544 27120 3596
rect 13544 3340 13596 3392
rect 13728 3340 13780 3392
rect 20444 3408 20496 3460
rect 24308 3476 24360 3528
rect 24768 3476 24820 3528
rect 25780 3451 25832 3460
rect 25780 3417 25789 3451
rect 25789 3417 25823 3451
rect 25823 3417 25832 3451
rect 25780 3408 25832 3417
rect 26516 3451 26568 3460
rect 26516 3417 26525 3451
rect 26525 3417 26559 3451
rect 26559 3417 26568 3451
rect 26516 3408 26568 3417
rect 16948 3383 17000 3392
rect 16948 3349 16957 3383
rect 16957 3349 16991 3383
rect 16991 3349 17000 3383
rect 16948 3340 17000 3349
rect 18236 3383 18288 3392
rect 18236 3349 18245 3383
rect 18245 3349 18279 3383
rect 18279 3349 18288 3383
rect 18236 3340 18288 3349
rect 18972 3340 19024 3392
rect 21180 3383 21232 3392
rect 21180 3349 21189 3383
rect 21189 3349 21223 3383
rect 21223 3349 21232 3383
rect 21180 3340 21232 3349
rect 23204 3340 23256 3392
rect 24124 3340 24176 3392
rect 5536 3238 5588 3290
rect 5600 3238 5652 3290
rect 5664 3238 5716 3290
rect 5728 3238 5780 3290
rect 14644 3238 14696 3290
rect 14708 3238 14760 3290
rect 14772 3238 14824 3290
rect 14836 3238 14888 3290
rect 23752 3238 23804 3290
rect 23816 3238 23868 3290
rect 23880 3238 23932 3290
rect 23944 3238 23996 3290
rect 4528 3136 4580 3188
rect 13728 3136 13780 3188
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 1492 3000 1544 3052
rect 480 2932 532 2984
rect 8668 3000 8720 3052
rect 9772 3068 9824 3120
rect 12256 3068 12308 3120
rect 12440 3068 12492 3120
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 3608 2975 3660 2984
rect 3608 2941 3617 2975
rect 3617 2941 3651 2975
rect 3651 2941 3660 2975
rect 3608 2932 3660 2941
rect 4160 2932 4212 2984
rect 6920 2975 6972 2984
rect 3240 2864 3292 2916
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 8300 2932 8352 2984
rect 10508 2932 10560 2984
rect 12348 3000 12400 3052
rect 12440 2932 12492 2984
rect 13544 2932 13596 2984
rect 13636 2932 13688 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 11980 2864 12032 2916
rect 12900 2864 12952 2916
rect 15936 2932 15988 2984
rect 18052 3136 18104 3188
rect 19156 3136 19208 3188
rect 24768 3136 24820 3188
rect 16396 3000 16448 3052
rect 17224 3000 17276 3052
rect 18420 3000 18472 3052
rect 19331 3043 19383 3052
rect 19331 3009 19349 3043
rect 19349 3009 19383 3043
rect 19331 3000 19383 3009
rect 16856 2932 16908 2984
rect 9588 2796 9640 2848
rect 12440 2796 12492 2848
rect 16028 2796 16080 2848
rect 18236 2864 18288 2916
rect 19892 2932 19944 2984
rect 20076 2932 20128 2984
rect 20720 2932 20772 2984
rect 22836 3000 22888 3052
rect 24124 2932 24176 2984
rect 25320 2932 25372 2984
rect 27344 2932 27396 2984
rect 20168 2864 20220 2916
rect 26240 2864 26292 2916
rect 17960 2796 18012 2848
rect 20352 2796 20404 2848
rect 20628 2796 20680 2848
rect 21640 2796 21692 2848
rect 23480 2796 23532 2848
rect 24768 2796 24820 2848
rect 26792 2839 26844 2848
rect 26792 2805 26801 2839
rect 26801 2805 26835 2839
rect 26835 2805 26844 2839
rect 26792 2796 26844 2805
rect 10090 2694 10142 2746
rect 10154 2694 10206 2746
rect 10218 2694 10270 2746
rect 10282 2694 10334 2746
rect 19198 2694 19250 2746
rect 19262 2694 19314 2746
rect 19326 2694 19378 2746
rect 19390 2694 19442 2746
rect 3608 2592 3660 2644
rect 4804 2524 4856 2576
rect 6460 2592 6512 2644
rect 9496 2592 9548 2644
rect 12532 2567 12584 2576
rect 12532 2533 12541 2567
rect 12541 2533 12575 2567
rect 12575 2533 12584 2567
rect 12532 2524 12584 2533
rect 12716 2592 12768 2644
rect 16764 2592 16816 2644
rect 16948 2524 17000 2576
rect 18420 2524 18472 2576
rect 19616 2524 19668 2576
rect 19984 2592 20036 2644
rect 20628 2592 20680 2644
rect 20168 2524 20220 2576
rect 21272 2592 21324 2644
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 2780 2456 2832 2508
rect 4620 2456 4672 2508
rect 5080 2456 5132 2508
rect 6000 2456 6052 2508
rect 6460 2456 6512 2508
rect 8024 2456 8076 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 9588 2499 9640 2508
rect 8484 2456 8536 2465
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 11520 2456 11572 2508
rect 11888 2456 11940 2508
rect 11244 2388 11296 2440
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 13820 2499 13872 2508
rect 12624 2456 12676 2465
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 14280 2456 14332 2508
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 17500 2456 17552 2508
rect 21180 2524 21232 2576
rect 23204 2567 23256 2576
rect 23204 2533 23213 2567
rect 23213 2533 23247 2567
rect 23247 2533 23256 2567
rect 23204 2524 23256 2533
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 7748 2320 7800 2372
rect 8300 2320 8352 2372
rect 9680 2320 9732 2372
rect 10600 2363 10652 2372
rect 10600 2329 10609 2363
rect 10609 2329 10643 2363
rect 10643 2329 10652 2363
rect 10600 2320 10652 2329
rect 15016 2320 15068 2372
rect 9772 2252 9824 2304
rect 13912 2295 13964 2304
rect 13912 2261 13921 2295
rect 13921 2261 13955 2295
rect 13955 2261 13964 2295
rect 13912 2252 13964 2261
rect 17132 2320 17184 2372
rect 20444 2456 20496 2508
rect 19984 2388 20036 2440
rect 23112 2499 23164 2508
rect 23112 2465 23121 2499
rect 23121 2465 23155 2499
rect 23155 2465 23164 2499
rect 23112 2456 23164 2465
rect 23388 2592 23440 2644
rect 24768 2592 24820 2644
rect 25872 2592 25924 2644
rect 24492 2524 24544 2576
rect 27068 2524 27120 2576
rect 23020 2388 23072 2440
rect 28540 2456 28592 2508
rect 20536 2320 20588 2372
rect 24952 2320 25004 2372
rect 28080 2320 28132 2372
rect 24124 2295 24176 2304
rect 24124 2261 24133 2295
rect 24133 2261 24167 2295
rect 24167 2261 24176 2295
rect 24124 2252 24176 2261
rect 5536 2150 5588 2202
rect 5600 2150 5652 2202
rect 5664 2150 5716 2202
rect 5728 2150 5780 2202
rect 14644 2150 14696 2202
rect 14708 2150 14760 2202
rect 14772 2150 14824 2202
rect 14836 2150 14888 2202
rect 23752 2150 23804 2202
rect 23816 2150 23868 2202
rect 23880 2150 23932 2202
rect 23944 2150 23996 2202
rect 11244 2048 11296 2100
rect 17684 2048 17736 2100
rect 4068 1980 4120 2032
rect 23112 1980 23164 2032
rect 8208 1912 8260 1964
rect 24124 1912 24176 1964
rect 1952 1844 2004 1896
rect 10508 1844 10560 1896
rect 13912 1844 13964 1896
rect 22192 1844 22244 1896
rect 7748 1776 7800 1828
rect 15016 1776 15068 1828
rect 21916 1776 21968 1828
rect 18696 1708 18748 1760
<< metal2 >>
rect 478 30924 534 31724
rect 938 30924 994 31724
rect 1858 30924 1914 31724
rect 2318 30924 2374 31724
rect 2778 30924 2834 31724
rect 3698 30924 3754 31724
rect 4158 30924 4214 31724
rect 5078 30924 5134 31724
rect 5538 30924 5594 31724
rect 5998 30924 6054 31724
rect 6918 30924 6974 31724
rect 7378 30924 7434 31724
rect 7838 30924 7894 31724
rect 8758 30924 8814 31724
rect 9218 30924 9274 31724
rect 9678 30924 9734 31724
rect 10598 30924 10654 31724
rect 11058 30924 11114 31724
rect 11518 30924 11574 31724
rect 12438 30924 12494 31724
rect 12898 30924 12954 31724
rect 13358 30924 13414 31724
rect 14278 30924 14334 31724
rect 14738 30924 14794 31724
rect 15198 30924 15254 31724
rect 16118 30924 16174 31724
rect 16578 30924 16634 31724
rect 17038 30924 17094 31724
rect 17958 30924 18014 31724
rect 18418 30924 18474 31724
rect 18878 30924 18934 31724
rect 19798 30924 19854 31724
rect 20258 30924 20314 31724
rect 20718 30924 20774 31724
rect 21638 30924 21694 31724
rect 22098 30924 22154 31724
rect 22558 30924 22614 31724
rect 23478 30924 23534 31724
rect 23938 30924 23994 31724
rect 24398 30924 24454 31724
rect 25318 30924 25374 31724
rect 25778 30924 25834 31724
rect 26238 30924 26294 31724
rect 27158 30924 27214 31724
rect 27618 30924 27674 31724
rect 28078 30924 28134 31724
rect 28998 30924 29054 31724
rect 492 28762 520 30924
rect 480 28756 532 28762
rect 480 28698 532 28704
rect 952 27606 980 30924
rect 1872 29458 1900 30924
rect 1872 29430 1992 29458
rect 1858 29336 1914 29345
rect 1858 29271 1914 29280
rect 1872 29102 1900 29271
rect 1964 29102 1992 29430
rect 1860 29096 1912 29102
rect 1860 29038 1912 29044
rect 1952 29096 2004 29102
rect 1952 29038 2004 29044
rect 2228 29028 2280 29034
rect 2228 28970 2280 28976
rect 2134 28656 2190 28665
rect 1768 28620 1820 28626
rect 2134 28591 2190 28600
rect 1768 28562 1820 28568
rect 1400 28008 1452 28014
rect 1398 27976 1400 27985
rect 1452 27976 1454 27985
rect 1398 27911 1454 27920
rect 940 27600 992 27606
rect 940 27542 992 27548
rect 1674 25936 1730 25945
rect 1674 25871 1676 25880
rect 1728 25871 1730 25880
rect 1676 25842 1728 25848
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1412 25265 1440 25298
rect 1398 25256 1454 25265
rect 1398 25191 1454 25200
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 17338 1440 17614
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1398 17096 1454 17105
rect 1398 17031 1454 17040
rect 1412 16658 1440 17031
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1412 14958 1440 14991
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1398 13016 1454 13025
rect 1398 12951 1454 12960
rect 1412 12782 1440 12951
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1412 9518 1440 9551
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 8945 1440 8978
rect 1398 8936 1454 8945
rect 1398 8871 1454 8880
rect 1504 8090 1532 24686
rect 1584 24676 1636 24682
rect 1584 24618 1636 24624
rect 1596 23662 1624 24618
rect 1676 24608 1728 24614
rect 1676 24550 1728 24556
rect 1688 23905 1716 24550
rect 1674 23896 1730 23905
rect 1674 23831 1730 23840
rect 1584 23656 1636 23662
rect 1584 23598 1636 23604
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 1688 20505 1716 21422
rect 1780 21298 1808 28562
rect 2148 28014 2176 28591
rect 2136 28008 2188 28014
rect 2136 27950 2188 27956
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 1950 26616 2006 26625
rect 1950 26551 1952 26560
rect 2004 26551 2006 26560
rect 1952 26522 2004 26528
rect 2148 26450 2176 26862
rect 2136 26444 2188 26450
rect 2136 26386 2188 26392
rect 2136 26240 2188 26246
rect 2240 26234 2268 28970
rect 2332 28762 2360 30924
rect 2412 29232 2464 29238
rect 2412 29174 2464 29180
rect 2320 28756 2372 28762
rect 2320 28698 2372 28704
rect 2240 26206 2360 26234
rect 2136 26182 2188 26188
rect 2148 25838 2176 26182
rect 2136 25832 2188 25838
rect 2136 25774 2188 25780
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 1860 23248 1912 23254
rect 1858 23216 1860 23225
rect 1912 23216 1914 23225
rect 1858 23151 1914 23160
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 22710 1992 22918
rect 1952 22704 2004 22710
rect 1952 22646 2004 22652
rect 2042 22536 2098 22545
rect 2042 22471 2044 22480
rect 2096 22471 2098 22480
rect 2044 22442 2096 22448
rect 2148 21486 2176 25094
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 1780 21270 2176 21298
rect 1950 21176 2006 21185
rect 1950 21111 1952 21120
rect 2004 21111 2006 21120
rect 1952 21082 2004 21088
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 1674 20496 1730 20505
rect 1674 20431 1730 20440
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1596 19310 1624 20334
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1596 18465 1624 18566
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17785 1624 18022
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1596 7954 1624 17478
rect 1688 11778 1716 19790
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1780 11880 1808 16730
rect 1872 16454 1900 20946
rect 1950 19816 2006 19825
rect 1950 19751 1952 19760
rect 2004 19751 2006 19760
rect 1952 19722 2004 19728
rect 2044 18148 2096 18154
rect 2044 18090 2096 18096
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 2056 16046 2084 18090
rect 2148 16250 2176 21270
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2240 19334 2268 19858
rect 2332 19514 2360 26206
rect 2424 23066 2452 29174
rect 2792 28150 2820 30924
rect 2870 30696 2926 30705
rect 2870 30631 2926 30640
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 2792 27606 2820 27950
rect 2780 27600 2832 27606
rect 2780 27542 2832 27548
rect 2884 27538 2912 30631
rect 3712 29306 3740 30924
rect 3700 29300 3752 29306
rect 3700 29242 3752 29248
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 2976 28150 3004 29106
rect 4172 28626 4200 30924
rect 5092 28626 5120 30924
rect 5552 30002 5580 30924
rect 5552 29974 5948 30002
rect 5510 29404 5806 29424
rect 5566 29402 5590 29404
rect 5646 29402 5670 29404
rect 5726 29402 5750 29404
rect 5588 29350 5590 29402
rect 5652 29350 5664 29402
rect 5726 29350 5728 29402
rect 5566 29348 5590 29350
rect 5646 29348 5670 29350
rect 5726 29348 5750 29350
rect 5510 29328 5806 29348
rect 5920 29238 5948 29974
rect 6012 29306 6040 30924
rect 6000 29300 6052 29306
rect 6000 29242 6052 29248
rect 5908 29232 5960 29238
rect 5908 29174 5960 29180
rect 5356 29028 5408 29034
rect 5356 28970 5408 28976
rect 5632 29028 5684 29034
rect 5632 28970 5684 28976
rect 3424 28620 3476 28626
rect 3424 28562 3476 28568
rect 4160 28620 4212 28626
rect 4160 28562 4212 28568
rect 5080 28620 5132 28626
rect 5080 28562 5132 28568
rect 2964 28144 3016 28150
rect 2964 28086 3016 28092
rect 2872 27532 2924 27538
rect 2872 27474 2924 27480
rect 2964 27328 3016 27334
rect 2964 27270 3016 27276
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2688 25288 2740 25294
rect 2688 25230 2740 25236
rect 2700 24818 2728 25230
rect 2884 24818 2912 25774
rect 2976 25430 3004 27270
rect 3332 25764 3384 25770
rect 3332 25706 3384 25712
rect 3344 25498 3372 25706
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 2964 25424 3016 25430
rect 2964 25366 3016 25372
rect 3148 25356 3200 25362
rect 3148 25298 3200 25304
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2516 23186 2544 24754
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 24342 2820 24550
rect 2884 24342 2912 24754
rect 3160 24750 3188 25298
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3160 24342 3188 24686
rect 3344 24682 3372 25298
rect 3332 24676 3384 24682
rect 3332 24618 3384 24624
rect 3344 24410 3372 24618
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 2780 24336 2832 24342
rect 2780 24278 2832 24284
rect 2872 24336 2924 24342
rect 2872 24278 2924 24284
rect 3148 24336 3200 24342
rect 3148 24278 3200 24284
rect 2884 23866 2912 24278
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 3056 23588 3108 23594
rect 3056 23530 3108 23536
rect 3068 23322 3096 23530
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 3160 23186 3188 24278
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 3148 23180 3200 23186
rect 3148 23122 3200 23128
rect 2424 23038 2544 23066
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2240 19306 2360 19334
rect 2332 18834 2360 19306
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 1858 14512 1914 14521
rect 1858 14447 1860 14456
rect 1912 14447 1914 14456
rect 1860 14418 1912 14424
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2042 14376 2098 14385
rect 1964 13870 1992 14350
rect 2042 14311 2044 14320
rect 2096 14311 2098 14320
rect 2044 14282 2096 14288
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 12220 1992 13806
rect 2240 13802 2268 15982
rect 2332 15706 2360 18770
rect 2424 16794 2452 19858
rect 2516 18630 2544 23038
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2240 13530 2268 13738
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12345 2084 12718
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2042 12336 2098 12345
rect 2042 12271 2098 12280
rect 1964 12192 2084 12220
rect 1780 11852 1900 11880
rect 1688 11750 1808 11778
rect 1674 11656 1730 11665
rect 1674 11591 1676 11600
rect 1728 11591 1730 11600
rect 1676 11562 1728 11568
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1688 9926 1716 10610
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9586 1716 9862
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1412 6905 1440 7890
rect 1596 7834 1624 7890
rect 1504 7806 1624 7834
rect 1504 7342 1532 7806
rect 1582 7576 1638 7585
rect 1582 7511 1584 7520
rect 1636 7511 1638 7520
rect 1584 7482 1636 7488
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1400 6248 1452 6254
rect 1398 6216 1400 6225
rect 1452 6216 1454 6225
rect 1398 6151 1454 6160
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4865 1440 5102
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1398 4856 1454 4865
rect 1596 4826 1624 4966
rect 1398 4791 1454 4800
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1780 4758 1808 11750
rect 1872 5574 1900 11852
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 10305 1992 10406
rect 1950 10296 2006 10305
rect 1950 10231 2006 10240
rect 2056 9042 2084 12192
rect 2240 11830 2268 12582
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2148 11354 2176 11630
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2148 10606 2176 11290
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8430 2084 8978
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2332 7342 2360 15302
rect 2412 14544 2464 14550
rect 2412 14486 2464 14492
rect 2424 13870 2452 14486
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2424 8974 2452 13806
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13462 2544 13670
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2424 8498 2452 8910
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2516 8430 2544 9318
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2424 6866 2452 7346
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6186 2176 6598
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 2148 5234 2176 6122
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2424 4758 2452 6802
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 940 3392 992 3398
rect 940 3334 992 3340
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 952 800 980 3334
rect 1412 800 1440 3878
rect 1780 3602 1808 4694
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2516 4282 2544 4626
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2608 3942 2636 23122
rect 3332 21412 3384 21418
rect 3332 21354 3384 21360
rect 3344 21146 3372 21354
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2700 19922 2728 20198
rect 2884 20058 2912 20266
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 3068 19990 3096 20878
rect 3056 19984 3108 19990
rect 3056 19926 3108 19932
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2872 18896 2924 18902
rect 2872 18838 2924 18844
rect 2884 18222 2912 18838
rect 3068 18222 3096 19246
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17134 2728 17478
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2792 16590 2820 17206
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2792 13190 2820 14894
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12850 2820 13126
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2792 12458 2820 12786
rect 2700 12430 2820 12458
rect 2700 12374 2728 12430
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2884 10266 2912 18158
rect 3068 17338 3096 18158
rect 3436 17882 3464 28562
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 4436 27872 4488 27878
rect 4436 27814 4488 27820
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4264 25498 4292 25638
rect 4252 25492 4304 25498
rect 4252 25434 4304 25440
rect 4344 25152 4396 25158
rect 4344 25094 4396 25100
rect 4356 24954 4384 25094
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4448 24274 4476 27814
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4540 24342 4568 24550
rect 4816 24410 4844 24618
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 4528 24336 4580 24342
rect 4528 24278 4580 24284
rect 4436 24268 4488 24274
rect 4436 24210 4488 24216
rect 4540 23662 4568 24278
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3896 23254 3924 23462
rect 3884 23248 3936 23254
rect 3884 23190 3936 23196
rect 3884 21616 3936 21622
rect 3884 21558 3936 21564
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3620 20398 3648 21422
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 16726 3004 16934
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 9178 2728 10066
rect 2884 9568 2912 10202
rect 2792 9540 2912 9568
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2792 9110 2820 9540
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2884 8634 2912 9386
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 6934 2728 7142
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2792 4554 2820 5034
rect 2884 4690 2912 7278
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2976 4570 3004 16662
rect 3160 16658 3188 17002
rect 3620 16794 3648 17070
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3804 16046 3832 21286
rect 3896 21010 3924 21558
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4250 21312 4306 21321
rect 4172 21078 4200 21286
rect 4250 21247 4306 21256
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 4264 20806 4292 21247
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3988 17270 4016 19858
rect 4264 18834 4292 20742
rect 4724 19281 4752 21558
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4908 21010 4936 21286
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4710 19272 4766 19281
rect 4710 19207 4766 19216
rect 4804 19236 4856 19242
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18902 4568 19110
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4724 18834 4752 19207
rect 4804 19178 4856 19184
rect 4816 18970 4844 19178
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4264 17762 4292 18770
rect 4264 17746 4384 17762
rect 4068 17740 4120 17746
rect 4264 17740 4396 17746
rect 4264 17734 4344 17740
rect 4068 17682 4120 17688
rect 4344 17682 4396 17688
rect 4080 17338 4108 17682
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4356 17270 4384 17682
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 3988 17134 4016 17206
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3896 16658 3924 17070
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 4356 16572 4384 17002
rect 4448 16726 4476 18770
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4540 17814 4568 18362
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4528 17808 4580 17814
rect 4528 17750 4580 17756
rect 4528 17672 4580 17678
rect 4632 17660 4660 18022
rect 4724 17746 4752 18770
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4816 17882 4844 18090
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4580 17632 4660 17660
rect 4528 17614 4580 17620
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4540 16572 4568 17614
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4632 16998 4660 17070
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4356 16544 4660 16572
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 14958 4200 15846
rect 4356 15162 4384 15914
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4356 14482 4384 15098
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3160 9654 3188 11630
rect 3252 11626 3280 13874
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 12782 4108 13670
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11694 3464 12038
rect 3712 11830 3740 12242
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3160 6662 3188 7210
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 5778 3188 6598
rect 3252 6458 3280 11562
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 10130 3556 10542
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9110 3648 9318
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3620 8362 3648 9046
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3436 6254 3464 6598
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2884 4542 3004 4570
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 2792 4078 2820 4111
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2884 4010 2912 4542
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 1504 3058 1532 3538
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1872 1465 1900 2450
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1964 1902 1992 2246
rect 1952 1896 2004 1902
rect 1952 1838 2004 1844
rect 1858 1456 1914 1465
rect 1858 1391 1914 1400
rect 2332 800 2360 3538
rect 2884 2990 2912 3946
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 800 2820 2450
rect 2976 2145 3004 4422
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3160 3505 3188 4014
rect 3146 3496 3202 3505
rect 3146 3431 3202 3440
rect 3620 2990 3648 8298
rect 3896 5370 3924 8366
rect 3988 7478 4016 12242
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11558 4108 11630
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 9586 4108 11494
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4172 8634 4200 13466
rect 4264 12986 4292 13738
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4356 11150 4384 13942
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4264 9518 4292 10406
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 9042 4292 9454
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4172 8378 4200 8570
rect 4080 8350 4200 8378
rect 4080 7546 4108 8350
rect 4356 7970 4384 11086
rect 4448 9450 4476 11154
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4540 9382 4568 10474
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4434 7984 4490 7993
rect 4356 7942 4434 7970
rect 4434 7919 4436 7928
rect 4488 7919 4490 7928
rect 4436 7890 4488 7896
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4080 7002 4108 7278
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4080 6458 4108 6938
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 6202 4200 7346
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4264 6730 4292 6802
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4264 6322 4292 6666
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4080 6186 4200 6202
rect 4068 6180 4200 6186
rect 4120 6174 4200 6180
rect 4068 6122 4120 6128
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3896 4758 3924 5306
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 4172 4622 4200 6174
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4264 4078 4292 6258
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 2962 2136 3018 2145
rect 2962 2071 3018 2080
rect 3252 800 3280 2858
rect 3620 2650 3648 2926
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 4080 2038 4108 3334
rect 4540 3194 4568 3946
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 4172 800 4200 2926
rect 4632 2774 4660 16544
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 4908 15366 4936 15914
rect 5000 15910 5028 28358
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5184 25294 5212 27406
rect 5264 25832 5316 25838
rect 5264 25774 5316 25780
rect 5276 25362 5304 25774
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5184 24818 5212 25230
rect 5276 24886 5304 25298
rect 5264 24880 5316 24886
rect 5264 24822 5316 24828
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 5184 24138 5212 24754
rect 5276 24206 5304 24822
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5172 24132 5224 24138
rect 5172 24074 5224 24080
rect 5184 22778 5212 24074
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5184 22098 5212 22714
rect 5276 22574 5304 23258
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5276 20602 5304 20946
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18426 5120 19246
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5368 17218 5396 28970
rect 5644 28762 5672 28970
rect 6932 28966 6960 30924
rect 6920 28960 6972 28966
rect 6920 28902 6972 28908
rect 5632 28756 5684 28762
rect 5632 28698 5684 28704
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 5510 28316 5806 28336
rect 5566 28314 5590 28316
rect 5646 28314 5670 28316
rect 5726 28314 5750 28316
rect 5588 28262 5590 28314
rect 5652 28262 5664 28314
rect 5726 28262 5728 28314
rect 5566 28260 5590 28262
rect 5646 28260 5670 28262
rect 5726 28260 5750 28262
rect 5510 28240 5806 28260
rect 6644 27872 6696 27878
rect 6644 27814 6696 27820
rect 5510 27228 5806 27248
rect 5566 27226 5590 27228
rect 5646 27226 5670 27228
rect 5726 27226 5750 27228
rect 5588 27174 5590 27226
rect 5652 27174 5664 27226
rect 5726 27174 5728 27226
rect 5566 27172 5590 27174
rect 5646 27172 5670 27174
rect 5726 27172 5750 27174
rect 5510 27152 5806 27172
rect 5510 26140 5806 26160
rect 5566 26138 5590 26140
rect 5646 26138 5670 26140
rect 5726 26138 5750 26140
rect 5588 26086 5590 26138
rect 5652 26086 5664 26138
rect 5726 26086 5728 26138
rect 5566 26084 5590 26086
rect 5646 26084 5670 26086
rect 5726 26084 5750 26086
rect 5510 26064 5806 26084
rect 5908 25832 5960 25838
rect 5908 25774 5960 25780
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5828 25430 5856 25638
rect 5816 25424 5868 25430
rect 5816 25366 5868 25372
rect 5510 25052 5806 25072
rect 5566 25050 5590 25052
rect 5646 25050 5670 25052
rect 5726 25050 5750 25052
rect 5588 24998 5590 25050
rect 5652 24998 5664 25050
rect 5726 24998 5728 25050
rect 5566 24996 5590 24998
rect 5646 24996 5670 24998
rect 5726 24996 5750 24998
rect 5510 24976 5806 24996
rect 5920 24342 5948 25774
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 5908 24336 5960 24342
rect 5908 24278 5960 24284
rect 5510 23964 5806 23984
rect 5566 23962 5590 23964
rect 5646 23962 5670 23964
rect 5726 23962 5750 23964
rect 5588 23910 5590 23962
rect 5652 23910 5664 23962
rect 5726 23910 5728 23962
rect 5566 23908 5590 23910
rect 5646 23908 5670 23910
rect 5726 23908 5750 23910
rect 5510 23888 5806 23908
rect 6000 23044 6052 23050
rect 6000 22986 6052 22992
rect 5510 22876 5806 22896
rect 5566 22874 5590 22876
rect 5646 22874 5670 22876
rect 5726 22874 5750 22876
rect 5588 22822 5590 22874
rect 5652 22822 5664 22874
rect 5726 22822 5728 22874
rect 5566 22820 5590 22822
rect 5646 22820 5670 22822
rect 5726 22820 5750 22822
rect 5510 22800 5806 22820
rect 5510 21788 5806 21808
rect 5566 21786 5590 21788
rect 5646 21786 5670 21788
rect 5726 21786 5750 21788
rect 5588 21734 5590 21786
rect 5652 21734 5664 21786
rect 5726 21734 5728 21786
rect 5566 21732 5590 21734
rect 5646 21732 5670 21734
rect 5726 21732 5750 21734
rect 5510 21712 5806 21732
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5736 21486 5764 21558
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5460 21321 5488 21422
rect 5446 21312 5502 21321
rect 5446 21247 5502 21256
rect 5828 21078 5856 21422
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 21078 5948 21286
rect 6012 21146 6040 22986
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 5816 21072 5868 21078
rect 5816 21014 5868 21020
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5816 20936 5868 20942
rect 5868 20884 5948 20890
rect 5816 20878 5948 20884
rect 5828 20862 5948 20878
rect 5510 20700 5806 20720
rect 5566 20698 5590 20700
rect 5646 20698 5670 20700
rect 5726 20698 5750 20700
rect 5588 20646 5590 20698
rect 5652 20646 5664 20698
rect 5726 20646 5728 20698
rect 5566 20644 5590 20646
rect 5646 20644 5670 20646
rect 5726 20644 5750 20646
rect 5510 20624 5806 20644
rect 5920 20602 5948 20862
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5552 19990 5580 20198
rect 5828 20058 5856 20266
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5540 19984 5592 19990
rect 5446 19952 5502 19961
rect 5540 19926 5592 19932
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5446 19887 5448 19896
rect 5500 19887 5502 19896
rect 5448 19858 5500 19864
rect 5510 19612 5806 19632
rect 5566 19610 5590 19612
rect 5646 19610 5670 19612
rect 5726 19610 5750 19612
rect 5588 19558 5590 19610
rect 5652 19558 5664 19610
rect 5726 19558 5728 19610
rect 5566 19556 5590 19558
rect 5646 19556 5670 19558
rect 5726 19556 5750 19558
rect 5510 19536 5806 19556
rect 5920 19310 5948 19926
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5510 18524 5806 18544
rect 5566 18522 5590 18524
rect 5646 18522 5670 18524
rect 5726 18522 5750 18524
rect 5588 18470 5590 18522
rect 5652 18470 5664 18522
rect 5726 18470 5728 18522
rect 5566 18468 5590 18470
rect 5646 18468 5670 18470
rect 5726 18468 5750 18470
rect 5510 18448 5806 18468
rect 6012 18222 6040 19858
rect 6104 18834 6132 25638
rect 6656 23186 6684 27814
rect 7116 26926 7144 28562
rect 7392 27606 7420 30924
rect 7852 29306 7880 30924
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 8772 29238 8800 30924
rect 8760 29232 8812 29238
rect 8760 29174 8812 29180
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7472 28688 7524 28694
rect 7470 28656 7472 28665
rect 7524 28656 7526 28665
rect 7470 28591 7526 28600
rect 7564 28620 7616 28626
rect 7564 28562 7616 28568
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7484 28014 7512 28358
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7576 27878 7604 28562
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 7380 27600 7432 27606
rect 7380 27542 7432 27548
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7564 27396 7616 27402
rect 7564 27338 7616 27344
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7392 26926 7420 27270
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7116 25362 7144 26862
rect 7392 25838 7420 26862
rect 7576 26858 7604 27338
rect 7668 27130 7696 27474
rect 7656 27124 7708 27130
rect 7656 27066 7708 27072
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 7484 25498 7512 25774
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 7380 25356 7432 25362
rect 7432 25316 7512 25344
rect 7380 25298 7432 25304
rect 7116 24886 7144 25298
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 7116 24274 7144 24822
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 7484 24070 7512 25316
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6092 18624 6144 18630
rect 6196 18612 6224 20742
rect 6288 20058 6316 22510
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6380 21146 6408 21422
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6380 19938 6408 21082
rect 6288 19910 6408 19938
rect 6288 19310 6316 19910
rect 6368 19848 6420 19854
rect 6472 19802 6500 22102
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 19990 6592 21830
rect 6656 21486 6684 22170
rect 6748 22094 6776 23462
rect 6932 22982 6960 23802
rect 7484 23662 7512 24006
rect 7576 23866 7604 24346
rect 7668 24342 7696 25094
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7564 23860 7616 23866
rect 7564 23802 7616 23808
rect 7576 23662 7604 23802
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 7576 22760 7604 23598
rect 7484 22732 7604 22760
rect 7208 22642 7420 22658
rect 7208 22636 7432 22642
rect 7208 22630 7380 22636
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22234 6868 22510
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6748 22066 6868 22094
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6748 21894 6776 21966
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6656 20466 6684 21422
rect 6748 21078 6776 21626
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6420 19796 6500 19802
rect 6368 19790 6500 19796
rect 6380 19774 6500 19790
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6144 18584 6224 18612
rect 6092 18566 6144 18572
rect 6104 18358 6132 18566
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5920 17814 5948 18022
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 6000 17536 6052 17542
rect 6104 17524 6132 18294
rect 6052 17496 6132 17524
rect 6000 17478 6052 17484
rect 5510 17436 5806 17456
rect 5566 17434 5590 17436
rect 5646 17434 5670 17436
rect 5726 17434 5750 17436
rect 5588 17382 5590 17434
rect 5652 17382 5664 17434
rect 5726 17382 5728 17434
rect 5566 17380 5590 17382
rect 5646 17380 5670 17382
rect 5726 17380 5750 17382
rect 5510 17360 5806 17380
rect 5276 17190 5396 17218
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15638 5212 15846
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4894 12744 4950 12753
rect 4894 12679 4950 12688
rect 4908 12306 4936 12679
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4724 11830 4752 12242
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 8634 4752 10542
rect 4816 10198 4844 10950
rect 4908 10742 4936 12242
rect 5000 12186 5028 13874
rect 5092 13530 5120 14214
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5092 13394 5120 13466
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12306 5120 13126
rect 5276 12434 5304 17190
rect 6012 16726 6040 17478
rect 6288 16794 6316 18906
rect 6380 18290 6408 19774
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 18698 6500 19246
rect 6748 18834 6776 19994
rect 6840 19310 6868 22066
rect 6932 21486 6960 22170
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6918 21312 6974 21321
rect 6918 21247 6974 21256
rect 6932 19922 6960 21247
rect 7024 19990 7052 22374
rect 7116 21690 7144 22442
rect 7208 22030 7236 22630
rect 7380 22578 7432 22584
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7300 22234 7328 22510
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7012 19984 7064 19990
rect 7012 19926 7064 19932
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 7116 19174 7144 20538
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5368 15910 5396 16662
rect 5510 16348 5806 16368
rect 5566 16346 5590 16348
rect 5646 16346 5670 16348
rect 5726 16346 5750 16348
rect 5588 16294 5590 16346
rect 5652 16294 5664 16346
rect 5726 16294 5728 16346
rect 5566 16292 5590 16294
rect 5646 16292 5670 16294
rect 5726 16292 5750 16294
rect 5510 16272 5806 16292
rect 6380 16182 6408 18226
rect 6472 16810 6500 18226
rect 6564 17338 6592 18770
rect 7024 18290 7052 19110
rect 7116 18766 7144 19110
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6472 16782 6592 16810
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6472 16182 6500 16662
rect 6368 16176 6420 16182
rect 6368 16118 6420 16124
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5828 15434 5856 15982
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5510 15260 5806 15280
rect 5566 15258 5590 15260
rect 5646 15258 5670 15260
rect 5726 15258 5750 15260
rect 5588 15206 5590 15258
rect 5652 15206 5664 15258
rect 5726 15206 5728 15258
rect 5566 15204 5590 15206
rect 5646 15204 5670 15206
rect 5726 15204 5750 15206
rect 5510 15184 5806 15204
rect 5920 14482 5948 15914
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 14006 5396 14214
rect 5510 14172 5806 14192
rect 5566 14170 5590 14172
rect 5646 14170 5670 14172
rect 5726 14170 5750 14172
rect 5588 14118 5590 14170
rect 5652 14118 5664 14170
rect 5726 14118 5728 14170
rect 5566 14116 5590 14118
rect 5646 14116 5670 14118
rect 5726 14116 5750 14118
rect 5510 14096 5806 14116
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5368 13870 5396 13942
rect 5552 13870 5580 13942
rect 5920 13938 5948 14418
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5552 13172 5580 13806
rect 6012 13734 6040 15642
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5920 13462 5948 13670
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5451 13144 5580 13172
rect 5451 12968 5479 13144
rect 5510 13084 5806 13104
rect 5566 13082 5590 13084
rect 5646 13082 5670 13084
rect 5726 13082 5750 13084
rect 5588 13030 5590 13082
rect 5652 13030 5664 13082
rect 5726 13030 5728 13082
rect 5566 13028 5590 13030
rect 5646 13028 5670 13030
rect 5726 13028 5750 13030
rect 5510 13008 5806 13028
rect 5451 12940 5488 12968
rect 5460 12782 5488 12940
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5184 12406 5304 12434
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5000 12158 5120 12186
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 5000 10674 5028 12038
rect 5092 11218 5120 12158
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4908 9178 4936 10542
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5000 9654 5028 10066
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5000 8906 5028 9590
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 5092 7954 5120 11154
rect 5184 8566 5212 12406
rect 5368 11626 5396 12718
rect 5736 12646 5764 12854
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5510 11996 5806 12016
rect 5566 11994 5590 11996
rect 5646 11994 5670 11996
rect 5726 11994 5750 11996
rect 5588 11942 5590 11994
rect 5652 11942 5664 11994
rect 5726 11942 5728 11994
rect 5566 11940 5590 11942
rect 5646 11940 5670 11942
rect 5726 11940 5750 11942
rect 5510 11920 5806 11940
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5276 9178 5304 10542
rect 5368 9518 5396 11562
rect 5920 11558 5948 12718
rect 6104 12646 6132 16050
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 6012 11354 6040 11630
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5510 10908 5806 10928
rect 5566 10906 5590 10908
rect 5646 10906 5670 10908
rect 5726 10906 5750 10908
rect 5588 10854 5590 10906
rect 5652 10854 5664 10906
rect 5726 10854 5728 10906
rect 5566 10852 5590 10854
rect 5646 10852 5670 10854
rect 5726 10852 5750 10854
rect 5510 10832 5806 10852
rect 5920 10266 5948 11154
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5510 9820 5806 9840
rect 5566 9818 5590 9820
rect 5646 9818 5670 9820
rect 5726 9818 5750 9820
rect 5588 9766 5590 9818
rect 5652 9766 5664 9818
rect 5726 9766 5728 9818
rect 5566 9764 5590 9766
rect 5646 9764 5670 9766
rect 5726 9764 5750 9766
rect 5510 9744 5806 9764
rect 5920 9722 5948 10066
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5368 9110 5396 9454
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5368 7970 5396 8842
rect 5552 8820 5580 9386
rect 6012 9042 6040 11290
rect 6104 10062 6132 11766
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5908 8832 5960 8838
rect 5552 8792 5908 8820
rect 5908 8774 5960 8780
rect 5510 8732 5806 8752
rect 5566 8730 5590 8732
rect 5646 8730 5670 8732
rect 5726 8730 5750 8732
rect 5588 8678 5590 8730
rect 5652 8678 5664 8730
rect 5726 8678 5728 8730
rect 5566 8676 5590 8678
rect 5646 8676 5670 8678
rect 5726 8676 5750 8678
rect 5510 8656 5806 8676
rect 5368 7954 5488 7970
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5368 7948 5500 7954
rect 5368 7942 5448 7948
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5000 7342 5028 7686
rect 5184 7342 5212 7822
rect 5368 7546 5396 7942
rect 5448 7890 5500 7896
rect 5510 7644 5806 7664
rect 5566 7642 5590 7644
rect 5646 7642 5670 7644
rect 5726 7642 5750 7644
rect 5588 7590 5590 7642
rect 5652 7590 5664 7642
rect 5726 7590 5728 7642
rect 5566 7588 5590 7590
rect 5646 7588 5670 7590
rect 5726 7588 5750 7590
rect 5510 7568 5806 7588
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5920 7410 5948 8774
rect 6090 7984 6146 7993
rect 6000 7948 6052 7954
rect 6090 7919 6092 7928
rect 6000 7890 6052 7896
rect 6144 7919 6146 7928
rect 6092 7890 6144 7896
rect 6012 7546 6040 7890
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6866 4752 7142
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4724 4078 4752 6802
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6390 5396 6734
rect 5510 6556 5806 6576
rect 5566 6554 5590 6556
rect 5646 6554 5670 6556
rect 5726 6554 5750 6556
rect 5588 6502 5590 6554
rect 5652 6502 5664 6554
rect 5726 6502 5728 6554
rect 5566 6500 5590 6502
rect 5646 6500 5670 6502
rect 5726 6500 5750 6502
rect 5510 6480 5806 6500
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5920 5914 5948 7210
rect 6196 6866 6224 15302
rect 6288 12170 6316 15642
rect 6472 15570 6500 16118
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6564 15348 6592 16782
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6656 15978 6684 16662
rect 6748 16114 6776 18158
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17882 6960 18090
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7116 17270 7144 18566
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6748 15638 6776 16050
rect 7024 15858 7052 16594
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7116 16046 7144 16458
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7104 15904 7156 15910
rect 7024 15852 7104 15858
rect 7024 15846 7156 15852
rect 7024 15830 7144 15846
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6472 15320 6592 15348
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6380 11830 6408 12718
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6361 6316 6598
rect 6274 6352 6330 6361
rect 6274 6287 6330 6296
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5510 5468 5806 5488
rect 5566 5466 5590 5468
rect 5646 5466 5670 5468
rect 5726 5466 5750 5468
rect 5588 5414 5590 5466
rect 5652 5414 5664 5466
rect 5726 5414 5728 5466
rect 5566 5412 5590 5414
rect 5646 5412 5670 5414
rect 5726 5412 5750 5414
rect 5510 5392 5806 5412
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4816 3602 4844 4558
rect 4908 4282 4936 4626
rect 6196 4486 6224 4626
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 5510 4380 5806 4400
rect 5566 4378 5590 4380
rect 5646 4378 5670 4380
rect 5726 4378 5750 4380
rect 5588 4326 5590 4378
rect 5652 4326 5664 4378
rect 5726 4326 5728 4378
rect 5566 4324 5590 4326
rect 5646 4324 5670 4326
rect 5726 4324 5750 4326
rect 5510 4304 5806 4324
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 6196 4146 6224 4422
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5368 3942 5396 4014
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5736 3738 5764 3878
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5920 3670 5948 3878
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5510 3292 5806 3312
rect 5566 3290 5590 3292
rect 5646 3290 5670 3292
rect 5726 3290 5750 3292
rect 5588 3238 5590 3290
rect 5652 3238 5664 3290
rect 5726 3238 5728 3290
rect 5566 3236 5590 3238
rect 5646 3236 5670 3238
rect 5726 3236 5750 3238
rect 5510 3216 5806 3236
rect 4632 2746 4844 2774
rect 4816 2582 4844 2746
rect 6472 2650 6500 15320
rect 6932 15026 6960 15506
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6656 13190 6684 13942
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6564 12306 6592 12854
rect 6656 12850 6684 13126
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6748 12646 6776 14282
rect 6840 13802 6868 14894
rect 6932 13802 6960 14962
rect 7116 14618 7144 15098
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7116 14074 7144 14554
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7208 13818 7236 21830
rect 7392 21486 7420 22374
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7484 21332 7512 22732
rect 7564 22568 7616 22574
rect 7564 22510 7616 22516
rect 7576 22098 7604 22510
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7300 21304 7512 21332
rect 7300 15638 7328 21304
rect 7576 20806 7604 21354
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7484 20058 7512 20266
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7380 19304 7432 19310
rect 7484 19281 7512 19858
rect 7576 19310 7604 20742
rect 7564 19304 7616 19310
rect 7380 19246 7432 19252
rect 7470 19272 7526 19281
rect 7392 18970 7420 19246
rect 7564 19246 7616 19252
rect 7470 19207 7526 19216
rect 7484 19122 7512 19207
rect 7484 19094 7604 19122
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18222 7420 18566
rect 7484 18222 7512 18906
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7392 17134 7420 18158
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7484 17066 7512 18158
rect 7576 17882 7604 19094
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7668 17218 7696 24142
rect 7576 17190 7696 17218
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 16946 7512 17002
rect 7392 16918 7512 16946
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 7116 13790 7236 13818
rect 6840 13530 6868 13738
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6656 9466 6684 12582
rect 6932 9568 6960 13262
rect 7116 13138 7144 13790
rect 7300 13258 7328 15574
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7116 13110 7328 13138
rect 7102 12880 7158 12889
rect 7102 12815 7158 12824
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10674 7052 11018
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6932 9540 7052 9568
rect 6564 9438 6684 9466
rect 6736 9444 6788 9450
rect 6564 7426 6592 9438
rect 6736 9386 6788 9392
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 9110 6684 9318
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6748 9042 6776 9386
rect 6932 9178 6960 9386
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6828 8424 6880 8430
rect 7024 8378 7052 9540
rect 6828 8366 6880 8372
rect 6840 7546 6868 8366
rect 6932 8350 7052 8378
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6564 7398 6684 7426
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6564 3398 6592 7278
rect 6656 6866 6684 7398
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6932 4826 6960 8350
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7342 7052 8230
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7116 7290 7144 12815
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7208 9178 7236 12650
rect 7300 12209 7328 13110
rect 7392 12238 7420 16918
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 13394 7512 14758
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7380 12232 7432 12238
rect 7286 12200 7342 12209
rect 7380 12174 7432 12180
rect 7286 12135 7342 12144
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11626 7328 12038
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7392 11150 7420 12174
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10606 7420 11086
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7484 9568 7512 13194
rect 7576 10062 7604 17190
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7668 14482 7696 15574
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13870 7696 14214
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7668 13190 7696 13330
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7300 9540 7512 9568
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7208 7410 7236 8978
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7116 7262 7236 7290
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6254 7052 6598
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7116 4010 7144 5102
rect 7208 4010 7236 7262
rect 7300 6730 7328 9540
rect 7484 9450 7512 9540
rect 7576 9518 7604 9862
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7392 7834 7420 9114
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7484 7954 7512 9046
rect 7576 8430 7604 9454
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7392 7806 7512 7834
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 6866 7420 7142
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7484 6662 7512 7806
rect 7668 7410 7696 13126
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 6934 7696 7346
rect 7760 6984 7788 28970
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8312 28626 8340 28902
rect 8574 28656 8630 28665
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 8300 28620 8352 28626
rect 8574 28591 8630 28600
rect 8300 28562 8352 28568
rect 7852 26926 7880 28562
rect 8588 28558 8616 28591
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 8760 27940 8812 27946
rect 8760 27882 8812 27888
rect 8668 27328 8720 27334
rect 8668 27270 8720 27276
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7852 25362 7880 26862
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 7840 25356 7892 25362
rect 7840 25298 7892 25304
rect 7852 24138 7880 25298
rect 8024 25288 8076 25294
rect 8024 25230 8076 25236
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7852 23730 7880 24074
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7852 19242 7880 19790
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7852 17218 7880 18294
rect 7944 18222 7972 20946
rect 8036 19334 8064 25230
rect 8220 25158 8248 25910
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 22658 8156 24550
rect 8220 22982 8248 25094
rect 8576 24676 8628 24682
rect 8576 24618 8628 24624
rect 8588 24410 8616 24618
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8128 22630 8248 22658
rect 8220 22094 8248 22630
rect 8128 22066 8248 22094
rect 8128 21894 8156 22066
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8220 19922 8248 21626
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8312 21010 8340 21354
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8312 20058 8340 20810
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8404 19922 8432 20742
rect 8496 19961 8524 21626
rect 8680 21010 8708 27270
rect 8772 27130 8800 27882
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 9232 26994 9260 30924
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9508 28626 9536 28902
rect 9692 28694 9720 30924
rect 9956 29572 10008 29578
rect 9956 29514 10008 29520
rect 9968 29102 9996 29514
rect 10612 29306 10640 30924
rect 10600 29300 10652 29306
rect 10600 29242 10652 29248
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 10968 29096 11020 29102
rect 10968 29038 11020 29044
rect 9864 29028 9916 29034
rect 9864 28970 9916 28976
rect 10692 29028 10744 29034
rect 10692 28970 10744 28976
rect 9680 28688 9732 28694
rect 9876 28665 9904 28970
rect 10064 28860 10360 28880
rect 10120 28858 10144 28860
rect 10200 28858 10224 28860
rect 10280 28858 10304 28860
rect 10142 28806 10144 28858
rect 10206 28806 10218 28858
rect 10280 28806 10282 28858
rect 10120 28804 10144 28806
rect 10200 28804 10224 28806
rect 10280 28804 10304 28806
rect 10064 28784 10360 28804
rect 9680 28630 9732 28636
rect 9862 28656 9918 28665
rect 9496 28620 9548 28626
rect 9862 28591 9918 28600
rect 10508 28620 10560 28626
rect 9496 28562 9548 28568
rect 10508 28562 10560 28568
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 9864 28484 9916 28490
rect 9864 28426 9916 28432
rect 9496 28008 9548 28014
rect 9496 27950 9548 27956
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9416 26926 9444 27406
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8956 24342 8984 24550
rect 8944 24336 8996 24342
rect 8944 24278 8996 24284
rect 8956 22574 8984 24278
rect 9416 23662 9444 26862
rect 9508 26586 9536 27950
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9692 26976 9720 27882
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9784 27538 9812 27814
rect 9876 27606 9904 28426
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9784 27169 9812 27474
rect 9770 27160 9826 27169
rect 9770 27095 9826 27104
rect 9864 27056 9916 27062
rect 9968 27044 9996 28494
rect 10244 28082 10272 28494
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10428 28150 10456 28358
rect 10416 28144 10468 28150
rect 10416 28086 10468 28092
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10416 27872 10468 27878
rect 10416 27814 10468 27820
rect 10064 27772 10360 27792
rect 10120 27770 10144 27772
rect 10200 27770 10224 27772
rect 10280 27770 10304 27772
rect 10142 27718 10144 27770
rect 10206 27718 10218 27770
rect 10280 27718 10282 27770
rect 10120 27716 10144 27718
rect 10200 27716 10224 27718
rect 10280 27716 10304 27718
rect 10064 27696 10360 27716
rect 10048 27056 10100 27062
rect 9968 27016 10048 27044
rect 9864 26998 9916 27004
rect 10048 26998 10100 27004
rect 9692 26948 9812 26976
rect 9678 26888 9734 26897
rect 9678 26823 9680 26832
rect 9732 26823 9734 26832
rect 9680 26794 9732 26800
rect 9588 26784 9640 26790
rect 9640 26732 9720 26738
rect 9588 26726 9720 26732
rect 9600 26710 9720 26726
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9508 26382 9536 26522
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9508 25838 9536 26318
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9508 24274 9536 25774
rect 9692 25498 9720 26710
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9692 23662 9720 24006
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9692 23186 9720 23598
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 8944 22568 8996 22574
rect 8944 22510 8996 22516
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8864 21486 8892 22374
rect 9140 22098 9168 22510
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9220 22432 9272 22438
rect 9220 22374 9272 22380
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8668 21004 8720 21010
rect 8668 20946 8720 20952
rect 8956 20806 8984 21558
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8588 19990 8616 20538
rect 8576 19984 8628 19990
rect 8482 19952 8538 19961
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 8392 19916 8444 19922
rect 8576 19926 8628 19932
rect 8482 19887 8538 19896
rect 8392 19858 8444 19864
rect 8036 19306 8156 19334
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7852 17190 7972 17218
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7852 16794 7880 17002
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7852 14634 7880 15914
rect 7944 14822 7972 17190
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7852 14606 7972 14634
rect 7840 14408 7892 14414
rect 7838 14376 7840 14385
rect 7892 14376 7894 14385
rect 7838 14311 7894 14320
rect 7852 12714 7880 14311
rect 7944 12889 7972 14606
rect 7930 12880 7986 12889
rect 7930 12815 7986 12824
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 8036 12442 8064 17070
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7838 12200 7894 12209
rect 7838 12135 7894 12144
rect 7852 9178 7880 12135
rect 8036 11830 8064 12378
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 8036 10674 8064 11766
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8128 10452 8156 19306
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18834 8432 19110
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8404 17882 8432 18634
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 11694 8248 17682
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 13530 8340 14894
rect 8588 14618 8616 15914
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8392 14612 8444 14618
rect 8576 14612 8628 14618
rect 8444 14572 8524 14600
rect 8392 14554 8444 14560
rect 8496 14074 8524 14572
rect 8576 14554 8628 14560
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8574 14376 8630 14385
rect 8574 14311 8576 14320
rect 8628 14311 8630 14320
rect 8576 14282 8628 14288
rect 8680 14278 8708 14554
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 12986 8340 13330
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8496 12782 8524 14010
rect 8772 12986 8800 14894
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8864 12866 8892 17138
rect 8956 15314 8984 20742
rect 9140 17338 9168 22034
rect 9232 21486 9260 22374
rect 9600 22098 9628 22442
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9692 21962 9720 22578
rect 9784 21962 9812 26948
rect 9876 26908 9904 26998
rect 10140 26920 10192 26926
rect 9876 26880 10140 26908
rect 10140 26862 10192 26868
rect 9860 26784 9912 26790
rect 9860 26726 9912 26732
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9876 26246 9904 26726
rect 9968 26518 9996 26726
rect 10064 26684 10360 26704
rect 10120 26682 10144 26684
rect 10200 26682 10224 26684
rect 10280 26682 10304 26684
rect 10142 26630 10144 26682
rect 10206 26630 10218 26682
rect 10280 26630 10282 26682
rect 10120 26628 10144 26630
rect 10200 26628 10224 26630
rect 10280 26628 10304 26630
rect 10064 26608 10360 26628
rect 9956 26512 10008 26518
rect 9956 26454 10008 26460
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9876 25362 9904 26182
rect 10428 25838 10456 27814
rect 10520 27674 10548 28562
rect 10704 28014 10732 28970
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 10508 27668 10560 27674
rect 10508 27610 10560 27616
rect 10980 27606 11008 29038
rect 11072 28694 11100 30924
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 11152 28416 11204 28422
rect 11072 28364 11152 28370
rect 11072 28358 11204 28364
rect 11072 28342 11192 28358
rect 10968 27600 11020 27606
rect 10506 27568 10562 27577
rect 10968 27542 11020 27548
rect 10506 27503 10508 27512
rect 10560 27503 10562 27512
rect 10508 27474 10560 27480
rect 10520 26858 10548 27474
rect 11072 27470 11100 28342
rect 11532 28014 11560 30924
rect 12452 29102 12480 30924
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 11520 28008 11572 28014
rect 11520 27950 11572 27956
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 10508 26852 10560 26858
rect 10508 26794 10560 26800
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 10064 25596 10360 25616
rect 10120 25594 10144 25596
rect 10200 25594 10224 25596
rect 10280 25594 10304 25596
rect 10142 25542 10144 25594
rect 10206 25542 10218 25594
rect 10280 25542 10282 25594
rect 10120 25540 10144 25542
rect 10200 25540 10224 25542
rect 10280 25540 10304 25542
rect 10064 25520 10360 25540
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 10060 24750 10088 25162
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10152 24750 10180 25094
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10064 24508 10360 24528
rect 10120 24506 10144 24508
rect 10200 24506 10224 24508
rect 10280 24506 10304 24508
rect 10142 24454 10144 24506
rect 10206 24454 10218 24506
rect 10280 24454 10282 24506
rect 10120 24452 10144 24454
rect 10200 24452 10224 24454
rect 10280 24452 10304 24454
rect 10064 24432 10360 24452
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9862 24168 9918 24177
rect 9862 24103 9918 24112
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9680 21616 9732 21622
rect 9678 21584 9680 21593
rect 9732 21584 9734 21593
rect 9678 21519 9734 21528
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9312 21344 9364 21350
rect 9312 21286 9364 21292
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9324 20398 9352 21286
rect 9416 21146 9444 21286
rect 9692 21146 9720 21422
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9496 21004 9548 21010
rect 9496 20946 9548 20952
rect 9508 20602 9536 20946
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9692 19174 9720 19994
rect 9784 19310 9812 21898
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9692 17218 9720 19110
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9784 17626 9812 18566
rect 9876 18426 9904 24103
rect 9968 23798 9996 24210
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 10520 23730 10548 26794
rect 11072 26450 11100 27406
rect 11900 26926 11928 27406
rect 11888 26920 11940 26926
rect 11888 26862 11940 26868
rect 11900 26518 11928 26862
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10888 25344 10916 25434
rect 10966 25392 11022 25401
rect 10888 25336 10966 25344
rect 10888 25316 10968 25336
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10612 24750 10640 25094
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10064 23420 10360 23440
rect 10120 23418 10144 23420
rect 10200 23418 10224 23420
rect 10280 23418 10304 23420
rect 10142 23366 10144 23418
rect 10206 23366 10218 23418
rect 10280 23366 10282 23418
rect 10120 23364 10144 23366
rect 10200 23364 10224 23366
rect 10280 23364 10304 23366
rect 10064 23344 10360 23364
rect 10428 23322 10456 23598
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 10232 22568 10284 22574
rect 9968 22528 10232 22556
rect 9968 22080 9996 22528
rect 10232 22510 10284 22516
rect 10064 22332 10360 22352
rect 10120 22330 10144 22332
rect 10200 22330 10224 22332
rect 10280 22330 10304 22332
rect 10142 22278 10144 22330
rect 10206 22278 10218 22330
rect 10280 22278 10282 22330
rect 10120 22276 10144 22278
rect 10200 22276 10224 22278
rect 10280 22276 10304 22278
rect 10064 22256 10360 22276
rect 10048 22092 10100 22098
rect 9968 22052 10048 22080
rect 10048 22034 10100 22040
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21486 9996 21830
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 10060 21332 10088 22034
rect 9968 21304 10088 21332
rect 9968 20040 9996 21304
rect 10064 21244 10360 21264
rect 10120 21242 10144 21244
rect 10200 21242 10224 21244
rect 10280 21242 10304 21244
rect 10142 21190 10144 21242
rect 10206 21190 10218 21242
rect 10280 21190 10282 21242
rect 10120 21188 10144 21190
rect 10200 21188 10224 21190
rect 10280 21188 10304 21190
rect 10064 21168 10360 21188
rect 10428 21078 10456 22714
rect 10520 21978 10548 22918
rect 10612 22778 10640 23598
rect 10704 23576 10732 24754
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10796 23730 10824 24618
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10784 23588 10836 23594
rect 10704 23548 10784 23576
rect 10784 23530 10836 23536
rect 10690 23216 10746 23225
rect 10690 23151 10746 23160
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10612 22098 10640 22442
rect 10704 22166 10732 23151
rect 10692 22160 10744 22166
rect 10692 22102 10744 22108
rect 10600 22092 10652 22098
rect 10600 22034 10652 22040
rect 10520 21950 10640 21978
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10520 20466 10548 21830
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10064 20156 10360 20176
rect 10120 20154 10144 20156
rect 10200 20154 10224 20156
rect 10280 20154 10304 20156
rect 10142 20102 10144 20154
rect 10206 20102 10218 20154
rect 10280 20102 10282 20154
rect 10120 20100 10144 20102
rect 10200 20100 10224 20102
rect 10280 20100 10304 20102
rect 10064 20080 10360 20100
rect 9968 20012 10088 20040
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 19514 9996 19858
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10060 19281 10088 20012
rect 10428 19922 10456 20334
rect 10508 20324 10560 20330
rect 10508 20266 10560 20272
rect 10520 20058 10548 20266
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10046 19272 10102 19281
rect 10046 19207 10102 19216
rect 10064 19068 10360 19088
rect 10120 19066 10144 19068
rect 10200 19066 10224 19068
rect 10280 19066 10304 19068
rect 10142 19014 10144 19066
rect 10206 19014 10218 19066
rect 10280 19014 10282 19066
rect 10120 19012 10144 19014
rect 10200 19012 10224 19014
rect 10280 19012 10304 19014
rect 10064 18992 10360 19012
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10244 18737 10272 18770
rect 10230 18728 10286 18737
rect 9956 18692 10008 18698
rect 10230 18663 10286 18672
rect 9956 18634 10008 18640
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9968 17746 9996 18634
rect 10336 18630 10364 18770
rect 10428 18698 10456 19858
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10064 17980 10360 18000
rect 10120 17978 10144 17980
rect 10200 17978 10224 17980
rect 10280 17978 10304 17980
rect 10142 17926 10144 17978
rect 10206 17926 10218 17978
rect 10280 17926 10282 17978
rect 10120 17924 10144 17926
rect 10200 17924 10224 17926
rect 10280 17924 10304 17926
rect 10064 17904 10360 17924
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9784 17598 9996 17626
rect 9862 17368 9918 17377
rect 9862 17303 9864 17312
rect 9916 17303 9918 17312
rect 9864 17274 9916 17280
rect 9600 17190 9720 17218
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 9048 15434 9076 17002
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 8956 15286 9076 15314
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8956 14278 8984 14826
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 9048 13258 9076 15286
rect 9600 15178 9628 17190
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9508 15150 9628 15178
rect 9508 15094 9536 15150
rect 9220 15088 9272 15094
rect 9220 15030 9272 15036
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9140 14929 9168 14962
rect 9126 14920 9182 14929
rect 9126 14855 9182 14864
rect 9126 14512 9182 14521
rect 9126 14447 9182 14456
rect 9140 14414 9168 14447
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8588 12838 8892 12866
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8588 12374 8616 12838
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8220 10742 8248 11290
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8128 10424 8248 10452
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8634 7880 8910
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7342 7880 7822
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7760 6956 7880 6984
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5302 7696 6190
rect 7760 5370 7788 6802
rect 7852 5914 7880 6956
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7116 3738 7144 3946
rect 7944 3942 7972 9998
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 4632 800 4660 2450
rect 5092 800 5120 2450
rect 5510 2204 5806 2224
rect 5566 2202 5590 2204
rect 5646 2202 5670 2204
rect 5726 2202 5750 2204
rect 5588 2150 5590 2202
rect 5652 2150 5664 2202
rect 5726 2150 5728 2202
rect 5566 2148 5590 2150
rect 5646 2148 5670 2150
rect 5726 2148 5750 2150
rect 5510 2128 5806 2148
rect 6012 800 6040 2450
rect 6472 800 6500 2450
rect 6932 800 6960 2926
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7760 1834 7788 2314
rect 7748 1828 7800 1834
rect 7748 1770 7800 1776
rect 7852 800 7880 3538
rect 8036 2990 8064 7142
rect 8128 6730 8156 7414
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8128 6458 8156 6666
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8036 2514 8064 2926
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8220 1970 8248 10424
rect 8312 10198 8340 11154
rect 8484 11008 8536 11014
rect 8482 10976 8484 10985
rect 8536 10976 8538 10985
rect 8482 10911 8538 10920
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8430 8524 8774
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8312 8090 8340 8366
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8312 5778 8340 8026
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 6186 8432 7346
rect 8482 6352 8538 6361
rect 8482 6287 8538 6296
rect 8496 6254 8524 6287
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8588 5817 8616 5850
rect 8574 5808 8630 5817
rect 8300 5772 8352 5778
rect 8574 5743 8630 5752
rect 8300 5714 8352 5720
rect 8312 5234 8340 5714
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4146 8340 5170
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8312 2990 8340 4082
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8496 2514 8524 4626
rect 8680 3534 8708 12718
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8772 11082 8800 11630
rect 9140 11150 9168 11698
rect 9036 11144 9088 11150
rect 9034 11112 9036 11121
rect 9128 11144 9180 11150
rect 9088 11112 9090 11121
rect 8760 11076 8812 11082
rect 9128 11086 9180 11092
rect 9034 11047 9090 11056
rect 8760 11018 8812 11024
rect 8772 10674 8800 11018
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 8362 8800 9318
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9140 8922 9168 9046
rect 9232 9042 9260 15030
rect 9692 14958 9720 17002
rect 9876 16998 9904 17274
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9784 15706 9812 16594
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9312 14952 9364 14958
rect 9680 14952 9732 14958
rect 9312 14894 9364 14900
rect 9586 14920 9642 14929
rect 9324 13530 9352 14894
rect 9680 14894 9732 14900
rect 9586 14855 9642 14864
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9416 9518 9444 14554
rect 9600 13462 9628 14855
rect 9692 14482 9720 14894
rect 9876 14618 9904 15846
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9968 14498 9996 17598
rect 10064 16892 10360 16912
rect 10120 16890 10144 16892
rect 10200 16890 10224 16892
rect 10280 16890 10304 16892
rect 10142 16838 10144 16890
rect 10206 16838 10218 16890
rect 10280 16838 10282 16890
rect 10120 16836 10144 16838
rect 10200 16836 10224 16838
rect 10280 16836 10304 16838
rect 10064 16816 10360 16836
rect 10064 15804 10360 15824
rect 10120 15802 10144 15804
rect 10200 15802 10224 15804
rect 10280 15802 10304 15804
rect 10142 15750 10144 15802
rect 10206 15750 10218 15802
rect 10280 15750 10282 15802
rect 10120 15748 10144 15750
rect 10200 15748 10224 15750
rect 10280 15748 10304 15750
rect 10064 15728 10360 15748
rect 10428 14890 10456 18634
rect 10508 18148 10560 18154
rect 10508 18090 10560 18096
rect 10520 17882 10548 18090
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10612 17762 10640 21950
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 10704 21690 10732 21898
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10796 21350 10824 23530
rect 10888 22982 10916 25316
rect 11020 25327 11022 25336
rect 10968 25298 11020 25304
rect 11072 24750 11100 26386
rect 11244 25900 11296 25906
rect 11244 25842 11296 25848
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 11164 25430 11192 25638
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 11256 25362 11284 25842
rect 11428 25764 11480 25770
rect 11428 25706 11480 25712
rect 11440 25498 11468 25706
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11900 25226 11928 26454
rect 12164 26240 12216 26246
rect 12164 26182 12216 26188
rect 12176 25838 12204 26182
rect 12072 25832 12124 25838
rect 12072 25774 12124 25780
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 12084 25294 12112 25774
rect 12268 25770 12296 27610
rect 12544 26874 12572 29242
rect 12912 29102 12940 30924
rect 12900 29096 12952 29102
rect 12900 29038 12952 29044
rect 12808 29028 12860 29034
rect 12808 28970 12860 28976
rect 12624 27532 12676 27538
rect 12624 27474 12676 27480
rect 12452 26846 12572 26874
rect 12348 26036 12400 26042
rect 12348 25978 12400 25984
rect 12256 25764 12308 25770
rect 12256 25706 12308 25712
rect 12268 25498 12296 25706
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 12084 24886 12112 25230
rect 12268 25158 12296 25298
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 11428 24880 11480 24886
rect 11428 24822 11480 24828
rect 12072 24880 12124 24886
rect 12072 24822 12124 24828
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10980 23322 11008 23598
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10888 21146 10916 22034
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10796 21026 10824 21082
rect 10980 21026 11008 23054
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 11072 22710 11100 22986
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10796 20998 11008 21026
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10704 19922 10732 20742
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10704 18578 10732 19450
rect 10796 19378 10824 20402
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10888 19174 10916 20998
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10704 18550 10824 18578
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10520 17734 10640 17762
rect 10704 17746 10732 18362
rect 10692 17740 10744 17746
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10064 14716 10360 14736
rect 10120 14714 10144 14716
rect 10200 14714 10224 14716
rect 10280 14714 10304 14716
rect 10142 14662 10144 14714
rect 10206 14662 10218 14714
rect 10280 14662 10282 14714
rect 10120 14660 10144 14662
rect 10200 14660 10224 14662
rect 10280 14660 10304 14662
rect 10064 14640 10360 14660
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9876 14470 9996 14498
rect 10416 14476 10468 14482
rect 9770 13832 9826 13841
rect 9770 13767 9826 13776
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9784 13394 9812 13767
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9876 12782 9904 14470
rect 10416 14418 10468 14424
rect 10322 14376 10378 14385
rect 10322 14311 10378 14320
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9864 12776 9916 12782
rect 9586 12744 9642 12753
rect 9642 12724 9864 12730
rect 9642 12718 9916 12724
rect 9642 12702 9904 12718
rect 9586 12679 9642 12688
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 11218 9720 12582
rect 9968 12306 9996 14214
rect 10336 13870 10364 14311
rect 10428 14278 10456 14418
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10064 13628 10360 13648
rect 10120 13626 10144 13628
rect 10200 13626 10224 13628
rect 10280 13626 10304 13628
rect 10142 13574 10144 13626
rect 10206 13574 10218 13626
rect 10280 13574 10282 13626
rect 10120 13572 10144 13574
rect 10200 13572 10224 13574
rect 10280 13572 10304 13574
rect 10064 13552 10360 13572
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10428 13258 10456 13330
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10520 13138 10548 17734
rect 10692 17682 10744 17688
rect 10796 17626 10824 18550
rect 10888 18222 10916 19110
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10888 17746 10916 18158
rect 10980 17882 11008 20470
rect 11072 20398 11100 22646
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 11164 21894 11192 22374
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19174 11100 19654
rect 11164 19310 11192 21830
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11256 19378 11284 20334
rect 11348 20058 11376 23666
rect 11440 22098 11468 24822
rect 12360 24721 12388 25978
rect 12346 24712 12402 24721
rect 12346 24647 12402 24656
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11624 19174 11652 22510
rect 11992 22234 12020 23122
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 12084 22574 12112 22918
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 12084 22166 12112 22510
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11716 21894 11744 21966
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 12268 20806 12296 22578
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12360 21486 12388 21626
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12360 20602 12388 21422
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11900 19281 11928 19858
rect 12256 19304 12308 19310
rect 11886 19272 11942 19281
rect 12256 19246 12308 19252
rect 11886 19207 11942 19216
rect 11980 19236 12032 19242
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10704 17598 10824 17626
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10876 17604 10928 17610
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10612 16794 10640 17274
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10704 15858 10732 17598
rect 10876 17546 10928 17552
rect 10888 16794 10916 17546
rect 10980 16794 11008 17614
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10612 15830 10732 15858
rect 10612 13841 10640 15830
rect 10692 15700 10744 15706
rect 10888 15688 10916 16730
rect 11072 16153 11100 19110
rect 11900 18834 11928 19207
rect 11980 19178 12032 19184
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11624 17814 11652 18090
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11900 17134 11928 18770
rect 11992 18630 12020 19178
rect 12268 18766 12296 19246
rect 12348 18896 12400 18902
rect 12346 18864 12348 18873
rect 12400 18864 12402 18873
rect 12346 18799 12402 18808
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16658 11560 17002
rect 12084 16726 12112 17682
rect 12268 17542 12296 18158
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12360 17202 12388 18090
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12360 16794 12388 17138
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11520 16652 11572 16658
rect 11440 16612 11520 16640
rect 11058 16144 11114 16153
rect 11058 16079 11114 16088
rect 10888 15660 11008 15688
rect 10692 15642 10744 15648
rect 10704 15502 10732 15642
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10692 15496 10744 15502
rect 10888 15473 10916 15506
rect 10980 15502 11008 15660
rect 10968 15496 11020 15502
rect 10692 15438 10744 15444
rect 10874 15464 10930 15473
rect 10704 15094 10732 15438
rect 10968 15438 11020 15444
rect 10874 15399 10876 15408
rect 10928 15399 10930 15408
rect 11060 15428 11112 15434
rect 10876 15370 10928 15376
rect 11060 15370 11112 15376
rect 10888 15339 10916 15370
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10782 14648 10838 14657
rect 11072 14618 11100 15370
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 10782 14583 10838 14592
rect 11060 14612 11112 14618
rect 10796 14414 10824 14583
rect 11060 14554 11112 14560
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13977 10824 14214
rect 10782 13968 10838 13977
rect 10782 13903 10838 13912
rect 10784 13864 10836 13870
rect 10598 13832 10654 13841
rect 10784 13806 10836 13812
rect 10598 13767 10654 13776
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10612 13394 10640 13466
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10428 13110 10548 13138
rect 10428 12918 10456 13110
rect 10612 13002 10640 13330
rect 10704 13326 10732 13738
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10520 12974 10640 13002
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10064 12540 10360 12560
rect 10120 12538 10144 12540
rect 10200 12538 10224 12540
rect 10280 12538 10304 12540
rect 10142 12486 10144 12538
rect 10206 12486 10218 12538
rect 10280 12486 10282 12538
rect 10120 12484 10144 12486
rect 10200 12484 10224 12486
rect 10280 12484 10304 12486
rect 10064 12464 10360 12484
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 10140 12300 10192 12306
rect 10520 12288 10548 12974
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10192 12260 10548 12288
rect 10140 12242 10192 12248
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11694 10364 12038
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10064 11452 10360 11472
rect 10120 11450 10144 11452
rect 10200 11450 10224 11452
rect 10280 11450 10304 11452
rect 10142 11398 10144 11450
rect 10206 11398 10218 11450
rect 10280 11398 10282 11450
rect 10120 11396 10144 11398
rect 10200 11396 10224 11398
rect 10280 11396 10304 11398
rect 10064 11376 10360 11396
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10130 9536 10950
rect 9968 10810 9996 11086
rect 10414 10976 10470 10985
rect 10414 10911 10470 10920
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9968 10690 9996 10746
rect 9876 10662 9996 10690
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9772 10124 9824 10130
rect 9876 10112 9904 10662
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 9968 10266 9996 10474
rect 10064 10364 10360 10384
rect 10120 10362 10144 10364
rect 10200 10362 10224 10364
rect 10280 10362 10304 10364
rect 10142 10310 10144 10362
rect 10206 10310 10218 10362
rect 10280 10310 10282 10362
rect 10120 10308 10144 10310
rect 10200 10308 10224 10310
rect 10280 10308 10304 10310
rect 10064 10288 10360 10308
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9824 10084 9904 10112
rect 9772 10066 9824 10072
rect 9692 10010 9720 10066
rect 9692 9982 9812 10010
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9140 8894 9260 8922
rect 9232 8566 9260 8894
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 9232 6254 9260 8502
rect 9416 8498 9444 9318
rect 9634 9104 9686 9110
rect 9784 9092 9812 9982
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9686 9064 9812 9092
rect 9634 9046 9686 9052
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9680 8424 9732 8430
rect 9784 8401 9812 9064
rect 9680 8366 9732 8372
rect 9770 8392 9826 8401
rect 9692 6798 9720 8366
rect 9770 8327 9826 8336
rect 9784 7018 9812 8327
rect 9968 7954 9996 9590
rect 10336 9489 10364 9930
rect 10322 9480 10378 9489
rect 10322 9415 10378 9424
rect 10064 9276 10360 9296
rect 10120 9274 10144 9276
rect 10200 9274 10224 9276
rect 10280 9274 10304 9276
rect 10142 9222 10144 9274
rect 10206 9222 10218 9274
rect 10280 9222 10282 9274
rect 10120 9220 10144 9222
rect 10200 9220 10224 9222
rect 10280 9220 10304 9222
rect 10064 9200 10360 9220
rect 10428 9178 10456 10911
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 8634 10088 8978
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10064 8188 10360 8208
rect 10120 8186 10144 8188
rect 10200 8186 10224 8188
rect 10280 8186 10304 8188
rect 10142 8134 10144 8186
rect 10206 8134 10218 8186
rect 10280 8134 10282 8186
rect 10120 8132 10144 8134
rect 10200 8132 10224 8134
rect 10280 8132 10304 8134
rect 10064 8112 10360 8132
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10064 7100 10360 7120
rect 10120 7098 10144 7100
rect 10200 7098 10224 7100
rect 10280 7098 10304 7100
rect 10142 7046 10144 7098
rect 10206 7046 10218 7098
rect 10280 7046 10282 7098
rect 10120 7044 10144 7046
rect 10200 7044 10224 7046
rect 10280 7044 10304 7046
rect 10064 7024 10360 7044
rect 9784 6990 9996 7018
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9140 4826 9168 6190
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5778 9536 6054
rect 9864 5908 9916 5914
rect 9784 5868 9864 5896
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9588 5704 9640 5710
rect 9784 5692 9812 5868
rect 9864 5850 9916 5856
rect 9862 5808 9918 5817
rect 9862 5743 9864 5752
rect 9916 5743 9918 5752
rect 9864 5714 9916 5720
rect 9968 5710 9996 6990
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6361 10180 6598
rect 10138 6352 10194 6361
rect 10138 6287 10194 6296
rect 10064 6012 10360 6032
rect 10120 6010 10144 6012
rect 10200 6010 10224 6012
rect 10280 6010 10304 6012
rect 10142 5958 10144 6010
rect 10206 5958 10218 6010
rect 10280 5958 10282 6010
rect 10120 5956 10144 5958
rect 10200 5956 10224 5958
rect 10280 5956 10304 5958
rect 10064 5936 10360 5956
rect 10428 5846 10456 8910
rect 10520 6798 10548 12260
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5914 10548 6190
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 9640 5664 9812 5692
rect 9956 5704 10008 5710
rect 9588 5646 9640 5652
rect 9956 5646 10008 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9508 4078 9536 5238
rect 9692 4758 9720 5510
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9784 4758 9812 5170
rect 10520 5098 10548 5714
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9588 3664 9640 3670
rect 9692 3641 9720 3946
rect 9588 3606 9640 3612
rect 9678 3632 9734 3641
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 3058 8708 3334
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8208 1964 8260 1970
rect 8208 1906 8260 1912
rect 8312 800 8340 2314
rect 8772 800 8800 3538
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9508 2650 9536 3402
rect 9600 2854 9628 3606
rect 9678 3567 9734 3576
rect 9784 3534 9812 4694
rect 9876 4690 9904 4966
rect 9968 4826 9996 5034
rect 10064 4924 10360 4944
rect 10120 4922 10144 4924
rect 10200 4922 10224 4924
rect 10280 4922 10304 4924
rect 10142 4870 10144 4922
rect 10206 4870 10218 4922
rect 10280 4870 10282 4922
rect 10120 4868 10144 4870
rect 10200 4868 10224 4870
rect 10280 4868 10304 4870
rect 10064 4848 10360 4868
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 10520 4282 10548 5034
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9876 3602 9904 3946
rect 10064 3836 10360 3856
rect 10120 3834 10144 3836
rect 10200 3834 10224 3836
rect 10280 3834 10304 3836
rect 10142 3782 10144 3834
rect 10206 3782 10218 3834
rect 10280 3782 10282 3834
rect 10120 3780 10144 3782
rect 10200 3780 10224 3782
rect 10280 3780 10304 3782
rect 10064 3760 10360 3780
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9692 3108 9720 3470
rect 9772 3120 9824 3126
rect 9692 3080 9772 3108
rect 9772 3062 9824 3068
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9600 2514 9628 2790
rect 10064 2748 10360 2768
rect 10120 2746 10144 2748
rect 10200 2746 10224 2748
rect 10280 2746 10304 2748
rect 10142 2694 10144 2746
rect 10206 2694 10218 2746
rect 10280 2694 10282 2746
rect 10120 2692 10144 2694
rect 10200 2692 10224 2694
rect 10280 2692 10304 2694
rect 10064 2672 10360 2692
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9770 2408 9826 2417
rect 9680 2372 9732 2378
rect 9770 2343 9826 2352
rect 9680 2314 9732 2320
rect 9692 800 9720 2314
rect 9784 2310 9812 2343
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 10428 1986 10456 4082
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10520 2990 10548 3334
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10612 2496 10640 12854
rect 10704 12442 10732 13262
rect 10796 13258 10824 13806
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10888 12782 10916 14486
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10980 13870 11008 14418
rect 11072 14006 11100 14554
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11164 14074 11192 14418
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12918 11008 13126
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10692 12436 10744 12442
rect 11072 12434 11100 13942
rect 11256 13852 11284 14350
rect 11348 14074 11376 14962
rect 11440 14890 11468 16612
rect 11520 16594 11572 16600
rect 12084 16046 12112 16662
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15502 12112 15982
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11336 13864 11388 13870
rect 11256 13824 11336 13852
rect 11256 13326 11284 13824
rect 11336 13806 11388 13812
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 10744 12406 10824 12434
rect 11072 12406 11284 12434
rect 10692 12378 10744 12384
rect 10796 12322 10824 12406
rect 10692 12300 10744 12306
rect 10796 12294 11008 12322
rect 10692 12242 10744 12248
rect 10704 11830 10732 12242
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10690 11112 10746 11121
rect 10690 11047 10746 11056
rect 10704 9518 10732 11047
rect 10796 10606 10824 12174
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10888 9654 10916 12174
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10796 8838 10824 9114
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8430 10824 8774
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 4826 10732 6734
rect 10796 6458 10824 8366
rect 10888 7546 10916 8978
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10980 7426 11008 12294
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 10674 11100 12038
rect 11256 11218 11284 12406
rect 11348 12374 11376 12922
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11348 11286 11376 11562
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11164 10810 11192 11154
rect 11440 11150 11468 14826
rect 11532 13802 11560 14962
rect 12162 13968 12218 13977
rect 12162 13903 12218 13912
rect 12176 13870 12204 13903
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11256 10062 11284 11018
rect 11348 10742 11376 11086
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11440 10538 11468 10950
rect 11428 10532 11480 10538
rect 11428 10474 11480 10480
rect 11440 10130 11468 10474
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11532 9874 11560 13738
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 11150 11652 13126
rect 12084 12918 12112 13806
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 11716 12442 11744 12854
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11992 11626 12020 12378
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11694 12112 12106
rect 12268 12102 12296 12854
rect 12452 12434 12480 26846
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12544 25430 12572 26726
rect 12636 26042 12664 27474
rect 12716 26852 12768 26858
rect 12716 26794 12768 26800
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12532 25424 12584 25430
rect 12532 25366 12584 25372
rect 12636 24886 12664 25638
rect 12728 25498 12756 26794
rect 12820 25514 12848 28970
rect 13372 28626 13400 30924
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 12992 28144 13044 28150
rect 12992 28086 13044 28092
rect 12716 25492 12768 25498
rect 12820 25486 12940 25514
rect 12716 25434 12768 25440
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12624 24880 12676 24886
rect 12624 24822 12676 24828
rect 12728 22574 12756 25230
rect 12820 25158 12848 25298
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22234 12756 22510
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12820 22094 12848 24074
rect 12728 22066 12848 22094
rect 12728 21486 12756 22066
rect 12820 21894 12848 22066
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12912 21554 12940 25486
rect 13004 24138 13032 28086
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 13096 27334 13124 27814
rect 14292 27606 14320 30924
rect 14752 30002 14780 30924
rect 14752 29974 15056 30002
rect 14618 29404 14914 29424
rect 14674 29402 14698 29404
rect 14754 29402 14778 29404
rect 14834 29402 14858 29404
rect 14696 29350 14698 29402
rect 14760 29350 14772 29402
rect 14834 29350 14836 29402
rect 14674 29348 14698 29350
rect 14754 29348 14778 29350
rect 14834 29348 14858 29350
rect 14618 29328 14914 29348
rect 15028 29102 15056 29974
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14372 28008 14424 28014
rect 14476 27962 14504 28494
rect 14618 28316 14914 28336
rect 14674 28314 14698 28316
rect 14754 28314 14778 28316
rect 14834 28314 14858 28316
rect 14696 28262 14698 28314
rect 14760 28262 14772 28314
rect 14834 28262 14836 28314
rect 14674 28260 14698 28262
rect 14754 28260 14778 28262
rect 14834 28260 14858 28262
rect 14618 28240 14914 28260
rect 15212 28014 15240 30924
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 14424 27956 14504 27962
rect 14372 27950 14504 27956
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 14384 27934 14504 27950
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 13360 27532 13412 27538
rect 13360 27474 13412 27480
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13280 26450 13308 27270
rect 13372 26926 13400 27474
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 13728 26512 13780 26518
rect 13728 26454 13780 26460
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13096 25294 13124 25434
rect 13188 25430 13216 26182
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13176 25424 13228 25430
rect 13176 25366 13228 25372
rect 13450 25392 13506 25401
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13004 23186 13032 23462
rect 13096 23186 13124 24686
rect 13188 24274 13216 25366
rect 13450 25327 13452 25336
rect 13504 25327 13506 25336
rect 13452 25298 13504 25304
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13176 23588 13228 23594
rect 13176 23530 13228 23536
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 12992 22092 13044 22098
rect 13096 22094 13124 23122
rect 13188 23100 13216 23530
rect 13280 23168 13308 24686
rect 13372 23730 13400 25230
rect 13648 24818 13676 25774
rect 13740 25498 13768 26454
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14004 25764 14056 25770
rect 14004 25706 14056 25712
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13740 25158 13768 25298
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13544 24676 13596 24682
rect 13544 24618 13596 24624
rect 13556 24410 13584 24618
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13740 23730 13768 25094
rect 13924 24886 13952 25434
rect 13912 24880 13964 24886
rect 13912 24822 13964 24828
rect 14016 24818 14044 25706
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 14108 24698 14136 25774
rect 14200 24750 14228 26726
rect 14280 25968 14332 25974
rect 14280 25910 14332 25916
rect 14292 25702 14320 25910
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14278 24848 14334 24857
rect 14278 24783 14334 24792
rect 14292 24750 14320 24783
rect 13924 24670 14136 24698
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 13924 24138 13952 24670
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13452 23180 13504 23186
rect 13280 23140 13452 23168
rect 13452 23122 13504 23128
rect 13188 23072 13308 23100
rect 13096 22066 13216 22094
rect 12992 22034 13044 22040
rect 13004 21894 13032 22034
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12636 21010 12664 21286
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13096 20058 13124 20334
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12544 17542 12572 18158
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12636 17814 12664 18022
rect 12624 17808 12676 17814
rect 12624 17750 12676 17756
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12544 16658 12572 17274
rect 12636 16726 12664 17614
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12728 16538 12756 19722
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 19446 13124 19654
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 13188 18873 13216 22066
rect 13280 22001 13308 23072
rect 13464 22234 13492 23122
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13266 21992 13322 22001
rect 13266 21927 13268 21936
rect 13320 21927 13322 21936
rect 13268 21898 13320 21904
rect 13280 21867 13308 21898
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13268 21344 13320 21350
rect 13266 21312 13268 21321
rect 13320 21312 13322 21321
rect 13266 21247 13322 21256
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13280 19786 13308 20470
rect 13372 19990 13400 20946
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13372 19174 13400 19926
rect 13464 19854 13492 21830
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13464 19446 13492 19790
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13268 18896 13320 18902
rect 13174 18864 13230 18873
rect 12992 18828 13044 18834
rect 13268 18838 13320 18844
rect 13174 18799 13230 18808
rect 12992 18770 13044 18776
rect 13004 18358 13032 18770
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13280 18154 13308 18838
rect 13372 18834 13400 19110
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13372 18290 13400 18770
rect 13556 18358 13584 22986
rect 13648 22506 13676 23462
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13636 22500 13688 22506
rect 13636 22442 13688 22448
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13648 20942 13676 21490
rect 13740 21486 13768 21830
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20942 13768 21286
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13648 18154 13676 20878
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13740 19922 13768 20266
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13740 19514 13768 19858
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13740 18698 13768 19450
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 18426 13768 18634
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12636 16510 12756 16538
rect 12636 15858 12664 16510
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 16046 12756 16390
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12636 15830 12756 15858
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12636 13530 12664 14894
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12452 12406 12572 12434
rect 12256 12096 12308 12102
rect 12308 12056 12388 12084
rect 12256 12038 12308 12044
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 9994 11652 11086
rect 11808 10130 11836 11154
rect 11992 10674 12020 11222
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 10985 12204 11018
rect 12162 10976 12218 10985
rect 12162 10911 12218 10920
rect 12360 10810 12388 12056
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 11980 10668 12032 10674
rect 12032 10628 12112 10656
rect 11980 10610 12032 10616
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9874 11744 9930
rect 11532 9846 11744 9874
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 9042 11100 9318
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11348 8634 11376 8978
rect 11624 8838 11652 8978
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10888 7398 11008 7426
rect 10888 6866 10916 7398
rect 11072 6866 11100 8298
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 6934 11192 7686
rect 11348 7002 11376 7890
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10888 5778 10916 6802
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 10888 5574 10916 5714
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 11440 5098 11468 5714
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11716 4729 11744 9846
rect 11808 7426 11836 10066
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11900 7546 11928 8978
rect 11992 8362 12020 10134
rect 12084 8430 12112 10628
rect 12360 10418 12388 10746
rect 12452 10538 12480 10950
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 12360 10390 12480 10418
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12176 9761 12204 10066
rect 12268 9994 12296 10066
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12162 9752 12218 9761
rect 12162 9687 12218 9696
rect 12176 9518 12204 9687
rect 12452 9586 12480 10390
rect 12544 10198 12572 12406
rect 12728 12170 12756 15830
rect 12820 15366 12848 16594
rect 12900 15632 12952 15638
rect 12900 15574 12952 15580
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12636 11218 12664 11562
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10470 12664 11154
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12544 9518 12572 9862
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12532 8424 12584 8430
rect 12636 8412 12664 10406
rect 12820 8922 12848 15302
rect 12912 11914 12940 15574
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13096 15065 13124 15098
rect 13082 15056 13138 15065
rect 13082 14991 13138 15000
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13734 13032 14214
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 12306 13032 13670
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12912 11886 13032 11914
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12912 11694 12940 11766
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11218 12940 11630
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 13004 11014 13032 11886
rect 13096 11558 13124 13874
rect 13188 11694 13216 15302
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12584 8384 12664 8412
rect 12728 8894 12848 8922
rect 12532 8366 12584 8372
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11808 7398 12020 7426
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 5778 11836 6734
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 4758 11836 5510
rect 11796 4752 11848 4758
rect 10690 4720 10746 4729
rect 10690 4655 10746 4664
rect 11702 4720 11758 4729
rect 11796 4694 11848 4700
rect 11702 4655 11758 4664
rect 10704 3602 10732 4655
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 11900 3516 11928 6666
rect 11992 4842 12020 7398
rect 12084 5166 12112 8366
rect 12176 8090 12204 8366
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12176 7342 12204 8026
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7342 12296 7686
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 6225 12296 6258
rect 12254 6216 12310 6225
rect 12254 6151 12310 6160
rect 12452 5710 12480 6802
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 5030 12112 5102
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11992 4814 12204 4842
rect 12176 4622 12204 4814
rect 12268 4758 12296 5034
rect 12452 4826 12480 5646
rect 12544 5302 12572 8366
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8022 12664 8230
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12636 5914 12664 6190
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12544 5166 12572 5238
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12176 4078 12204 4558
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 11980 3528 12032 3534
rect 11900 3488 11980 3516
rect 11900 2514 11928 3488
rect 11980 3470 12032 3476
rect 12254 3224 12310 3233
rect 12254 3159 12310 3168
rect 12268 3126 12296 3159
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12360 3058 12388 3975
rect 12452 3670 12480 4218
rect 12530 4176 12586 4185
rect 12530 4111 12586 4120
rect 12544 4010 12572 4111
rect 12636 4078 12664 4966
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12728 3890 12756 8894
rect 12912 8838 12940 8978
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12820 7478 12848 8774
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12912 6254 12940 8774
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12820 5896 12848 6190
rect 12900 5908 12952 5914
rect 12820 5868 12900 5896
rect 12900 5850 12952 5856
rect 13004 5778 13032 6598
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13096 5166 13124 7890
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12820 4690 12848 5102
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12820 4282 12848 4626
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12992 3936 13044 3942
rect 12636 3862 12848 3890
rect 12992 3878 13044 3884
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12452 3126 12480 3606
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12440 2984 12492 2990
rect 12438 2952 12440 2961
rect 12492 2952 12494 2961
rect 11980 2916 12032 2922
rect 12438 2887 12494 2896
rect 11980 2858 12032 2864
rect 10152 1958 10456 1986
rect 10520 2468 10640 2496
rect 11520 2508 11572 2514
rect 10152 800 10180 1958
rect 10520 1902 10548 2468
rect 11520 2450 11572 2456
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10612 800 10640 2314
rect 11256 2106 11284 2382
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 11532 800 11560 2450
rect 11992 800 12020 2858
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 800 12480 2790
rect 12544 2582 12572 3402
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12636 2514 12664 3862
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12728 2650 12756 3538
rect 12820 3346 12848 3862
rect 13004 3777 13032 3878
rect 12990 3768 13046 3777
rect 12900 3732 12952 3738
rect 12990 3703 13046 3712
rect 12900 3674 12952 3680
rect 12912 3641 12940 3674
rect 12898 3632 12954 3641
rect 13096 3618 13124 4082
rect 13188 4049 13216 11018
rect 13280 7562 13308 17478
rect 13372 15892 13400 18090
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13464 16182 13492 16662
rect 13556 16658 13584 16934
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13464 16046 13492 16118
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13372 15864 13492 15892
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13372 15162 13400 15506
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13464 14482 13492 15864
rect 13648 14634 13676 16934
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15570 13768 15846
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13832 15366 13860 22646
rect 13924 19310 13952 24074
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13924 17746 13952 18770
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13556 14606 13676 14634
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13464 14006 13492 14282
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13464 12782 13492 13942
rect 13556 12918 13584 14606
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13556 12434 13584 12854
rect 13464 12406 13584 12434
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11762 13400 12038
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13464 11694 13492 12406
rect 13452 11688 13504 11694
rect 13372 11636 13452 11642
rect 13372 11630 13504 11636
rect 13372 11614 13492 11630
rect 13372 10690 13400 11614
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11354 13584 11494
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13464 10810 13492 11222
rect 13648 11082 13676 14418
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13190 13768 14214
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13832 12374 13860 15302
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13924 12986 13952 13806
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14016 12442 14044 24006
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 14108 22778 14136 23598
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14200 23186 14228 23462
rect 14292 23304 14320 24686
rect 14384 24342 14412 27406
rect 14476 26450 14504 27934
rect 15292 27940 15344 27946
rect 15292 27882 15344 27888
rect 15304 27674 15332 27882
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15108 27668 15160 27674
rect 15292 27668 15344 27674
rect 15160 27628 15240 27656
rect 15108 27610 15160 27616
rect 15106 27568 15162 27577
rect 15212 27538 15240 27628
rect 15292 27610 15344 27616
rect 15396 27606 15424 27814
rect 15580 27606 15608 29650
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15568 27600 15620 27606
rect 15568 27542 15620 27548
rect 15028 27512 15106 27520
rect 15028 27492 15108 27512
rect 14618 27228 14914 27248
rect 14674 27226 14698 27228
rect 14754 27226 14778 27228
rect 14834 27226 14858 27228
rect 14696 27174 14698 27226
rect 14760 27174 14772 27226
rect 14834 27174 14836 27226
rect 14674 27172 14698 27174
rect 14754 27172 14778 27174
rect 14834 27172 14858 27174
rect 14618 27152 14914 27172
rect 14464 26444 14516 26450
rect 14464 26386 14516 26392
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14476 25906 14504 26250
rect 14618 26140 14914 26160
rect 14674 26138 14698 26140
rect 14754 26138 14778 26140
rect 14834 26138 14858 26140
rect 14696 26086 14698 26138
rect 14760 26086 14772 26138
rect 14834 26086 14836 26138
rect 14674 26084 14698 26086
rect 14754 26084 14778 26086
rect 14834 26084 14858 26086
rect 14618 26064 14914 26084
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14618 25052 14914 25072
rect 14674 25050 14698 25052
rect 14754 25050 14778 25052
rect 14834 25050 14858 25052
rect 14696 24998 14698 25050
rect 14760 24998 14772 25050
rect 14834 24998 14836 25050
rect 14674 24996 14698 24998
rect 14754 24996 14778 24998
rect 14834 24996 14858 24998
rect 14618 24976 14914 24996
rect 14924 24880 14976 24886
rect 14922 24848 14924 24857
rect 14976 24848 14978 24857
rect 14922 24783 14978 24792
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14618 23964 14914 23984
rect 14674 23962 14698 23964
rect 14754 23962 14778 23964
rect 14834 23962 14858 23964
rect 14696 23910 14698 23962
rect 14760 23910 14772 23962
rect 14834 23910 14836 23962
rect 14674 23908 14698 23910
rect 14754 23908 14778 23910
rect 14834 23908 14858 23910
rect 14618 23888 14914 23908
rect 15028 23526 15056 27492
rect 15160 27503 15162 27512
rect 15200 27532 15252 27538
rect 15108 27474 15160 27480
rect 15200 27474 15252 27480
rect 15580 26994 15608 27542
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15120 25158 15148 26862
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15120 24188 15148 25094
rect 15212 24410 15240 25366
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15304 24206 15332 24686
rect 15488 24274 15516 26862
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15580 26518 15608 26726
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15672 24954 15700 25774
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15200 24200 15252 24206
rect 15120 24160 15200 24188
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 14462 23352 14518 23361
rect 14292 23276 14412 23304
rect 15120 23322 15148 24160
rect 15200 24142 15252 24148
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15488 23730 15516 24210
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 14462 23287 14518 23296
rect 15108 23316 15160 23322
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14094 21312 14150 21321
rect 14094 21247 14150 21256
rect 14108 20466 14136 21247
rect 14200 20806 14228 21422
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14108 19378 14136 19722
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14108 18970 14136 19314
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14200 18086 14228 20538
rect 14292 20262 14320 21286
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17649 14228 18022
rect 14292 17746 14320 20198
rect 14384 17814 14412 23276
rect 14476 23254 14504 23287
rect 15108 23258 15160 23264
rect 14464 23248 14516 23254
rect 14464 23190 14516 23196
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14844 23089 14872 23122
rect 15016 23112 15068 23118
rect 14830 23080 14886 23089
rect 15016 23054 15068 23060
rect 14830 23015 14886 23024
rect 14618 22876 14914 22896
rect 14674 22874 14698 22876
rect 14754 22874 14778 22876
rect 14834 22874 14858 22876
rect 14696 22822 14698 22874
rect 14760 22822 14772 22874
rect 14834 22822 14836 22874
rect 14674 22820 14698 22822
rect 14754 22820 14778 22822
rect 14834 22820 14858 22822
rect 14618 22800 14914 22820
rect 15028 22778 15056 23054
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 15212 21894 15240 23598
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15304 22098 15332 23530
rect 15488 22710 15516 23666
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15292 22092 15344 22098
rect 15488 22094 15516 22510
rect 15292 22034 15344 22040
rect 15396 22066 15516 22094
rect 15304 21894 15332 22034
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 14618 21788 14914 21808
rect 14674 21786 14698 21788
rect 14754 21786 14778 21788
rect 14834 21786 14858 21788
rect 14696 21734 14698 21786
rect 14760 21734 14772 21786
rect 14834 21734 14836 21786
rect 14674 21732 14698 21734
rect 14754 21732 14778 21734
rect 14834 21732 14858 21734
rect 14618 21712 14914 21732
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14844 21010 14872 21558
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14476 19514 14504 20946
rect 14844 20874 14872 20946
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14618 20700 14914 20720
rect 14674 20698 14698 20700
rect 14754 20698 14778 20700
rect 14834 20698 14858 20700
rect 14696 20646 14698 20698
rect 14760 20646 14772 20698
rect 14834 20646 14836 20698
rect 14674 20644 14698 20646
rect 14754 20644 14778 20646
rect 14834 20644 14858 20646
rect 14618 20624 14914 20644
rect 15028 19786 15056 21490
rect 15212 21350 15240 21830
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15120 21162 15148 21286
rect 15120 21134 15240 21162
rect 15212 21010 15240 21134
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 15120 20602 15148 20878
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15304 20398 15332 21422
rect 15396 21026 15424 22066
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15488 21486 15516 21830
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15396 21010 15516 21026
rect 15396 21004 15528 21010
rect 15396 20998 15476 21004
rect 15476 20946 15528 20952
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15488 20754 15516 20946
rect 15580 20874 15608 24754
rect 15660 24744 15712 24750
rect 15658 24712 15660 24721
rect 15712 24712 15714 24721
rect 15658 24647 15714 24656
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 14618 19612 14914 19632
rect 14674 19610 14698 19612
rect 14754 19610 14778 19612
rect 14834 19610 14858 19612
rect 14696 19558 14698 19610
rect 14760 19558 14772 19610
rect 14834 19558 14836 19610
rect 14674 19556 14698 19558
rect 14754 19556 14778 19558
rect 14834 19556 14858 19558
rect 14618 19536 14914 19556
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14476 19334 14504 19450
rect 14476 19306 14688 19334
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18873 14504 19110
rect 14660 18873 14688 19306
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14462 18864 14518 18873
rect 14462 18799 14518 18808
rect 14646 18864 14702 18873
rect 14752 18834 14780 19178
rect 15028 18834 15056 19722
rect 15120 19530 15148 20334
rect 15304 19922 15332 20334
rect 15396 20058 15424 20742
rect 15488 20726 15608 20754
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15120 19502 15240 19530
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 14646 18799 14702 18808
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14476 18290 14504 18702
rect 14618 18524 14914 18544
rect 14674 18522 14698 18524
rect 14754 18522 14778 18524
rect 14834 18522 14858 18524
rect 14696 18470 14698 18522
rect 14760 18470 14772 18522
rect 14834 18470 14836 18522
rect 14674 18468 14698 18470
rect 14754 18468 14778 18470
rect 14834 18468 14858 18470
rect 14618 18448 14914 18468
rect 15028 18358 15056 18770
rect 15120 18766 15148 19314
rect 15212 19310 15240 19502
rect 15200 19304 15252 19310
rect 15488 19281 15516 19790
rect 15200 19246 15252 19252
rect 15474 19272 15530 19281
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15212 18630 15240 19246
rect 15474 19207 15530 19216
rect 15290 18728 15346 18737
rect 15290 18663 15346 18672
rect 15200 18624 15252 18630
rect 15120 18572 15200 18578
rect 15120 18566 15252 18572
rect 15120 18550 15240 18566
rect 15016 18352 15068 18358
rect 15016 18294 15068 18300
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14186 17640 14242 17649
rect 14186 17575 14242 17584
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14108 16969 14136 17478
rect 14200 17066 14228 17575
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14094 16960 14150 16969
rect 14094 16895 14150 16904
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14929 14136 14962
rect 14200 14958 14228 15370
rect 14188 14952 14240 14958
rect 14094 14920 14150 14929
rect 14188 14894 14240 14900
rect 14094 14855 14150 14864
rect 14186 14512 14242 14521
rect 14186 14447 14242 14456
rect 14200 14006 14228 14447
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14108 12646 14136 12922
rect 14200 12714 14228 13942
rect 14292 13802 14320 17682
rect 14384 15638 14412 17750
rect 15028 17610 15056 18294
rect 15120 18222 15148 18550
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14464 17536 14516 17542
rect 15200 17536 15252 17542
rect 14464 17478 14516 17484
rect 15120 17496 15200 17524
rect 14476 16658 14504 17478
rect 14618 17436 14914 17456
rect 14674 17434 14698 17436
rect 14754 17434 14778 17436
rect 14834 17434 14858 17436
rect 14696 17382 14698 17434
rect 14760 17382 14772 17434
rect 14834 17382 14836 17434
rect 14674 17380 14698 17382
rect 14754 17380 14778 17382
rect 14834 17380 14858 17382
rect 14618 17360 14914 17380
rect 15120 16658 15148 17496
rect 15200 17478 15252 17484
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14476 15450 14504 16594
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14618 16348 14914 16368
rect 14674 16346 14698 16348
rect 14754 16346 14778 16348
rect 14834 16346 14858 16348
rect 14696 16294 14698 16346
rect 14760 16294 14772 16346
rect 14834 16294 14836 16346
rect 14674 16292 14698 16294
rect 14754 16292 14778 16294
rect 14834 16292 14858 16294
rect 14618 16272 14914 16292
rect 15028 15978 15056 16526
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14384 15422 14504 15450
rect 14384 13870 14412 15422
rect 14618 15260 14914 15280
rect 14674 15258 14698 15260
rect 14754 15258 14778 15260
rect 14834 15258 14858 15260
rect 14696 15206 14698 15258
rect 14760 15206 14772 15258
rect 14834 15206 14836 15258
rect 14674 15204 14698 15206
rect 14754 15204 14778 15206
rect 14834 15204 14858 15206
rect 14618 15184 14914 15204
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14476 14822 14504 15098
rect 14740 14952 14792 14958
rect 14924 14952 14976 14958
rect 14740 14894 14792 14900
rect 14830 14920 14886 14929
rect 14752 14822 14780 14894
rect 15028 14940 15056 15914
rect 14976 14912 15056 14940
rect 14924 14894 14976 14900
rect 14830 14855 14832 14864
rect 14884 14855 14886 14864
rect 14832 14826 14884 14832
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14922 14784 14978 14793
rect 14752 14482 14780 14758
rect 14922 14719 14978 14728
rect 14936 14482 14964 14719
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 14464 14408 14516 14414
rect 14752 14385 14780 14418
rect 14464 14350 14516 14356
rect 14738 14376 14794 14385
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14476 13802 14504 14350
rect 14738 14311 14794 14320
rect 14618 14172 14914 14192
rect 14674 14170 14698 14172
rect 14754 14170 14778 14172
rect 14834 14170 14858 14172
rect 14696 14118 14698 14170
rect 14760 14118 14772 14170
rect 14834 14118 14836 14170
rect 14674 14116 14698 14118
rect 14754 14116 14778 14118
rect 14834 14116 14858 14118
rect 14618 14096 14914 14116
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14292 12782 14320 13738
rect 14618 13084 14914 13104
rect 14674 13082 14698 13084
rect 14754 13082 14778 13084
rect 14834 13082 14858 13084
rect 14696 13030 14698 13082
rect 14760 13030 14772 13082
rect 14834 13030 14836 13082
rect 14674 13028 14698 13030
rect 14754 13028 14778 13030
rect 14834 13028 14858 13030
rect 14618 13008 14914 13028
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 14108 11626 14136 12582
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13372 10662 13492 10690
rect 13464 9586 13492 10662
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13464 9042 13492 9522
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13556 8401 13584 10406
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13648 8974 13676 9386
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9178 13768 9318
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8430 13676 8910
rect 13636 8424 13688 8430
rect 13542 8392 13598 8401
rect 13636 8366 13688 8372
rect 13542 8327 13544 8336
rect 13596 8327 13598 8336
rect 13544 8298 13596 8304
rect 13648 8294 13676 8366
rect 13648 8266 13768 8294
rect 13280 7534 13676 7562
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13280 5710 13308 7414
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13266 4720 13322 4729
rect 13266 4655 13268 4664
rect 13320 4655 13322 4664
rect 13268 4626 13320 4632
rect 13372 4214 13400 7346
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13464 4826 13492 5034
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13556 4282 13584 4966
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13004 3602 13124 3618
rect 12898 3567 12954 3576
rect 12992 3596 13124 3602
rect 13044 3590 13124 3596
rect 12992 3538 13044 3544
rect 13188 3466 13216 3878
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 13280 3346 13308 3538
rect 12820 3318 13308 3346
rect 12898 3224 12954 3233
rect 12898 3159 12954 3168
rect 12912 2922 12940 3159
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13372 800 13400 3946
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13556 2990 13584 3334
rect 13648 2990 13676 7534
rect 13740 6186 13768 8266
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13832 5846 13860 11562
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13924 9761 13952 10746
rect 13910 9752 13966 9761
rect 13910 9687 13966 9696
rect 13924 9654 13952 9687
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14200 8537 14228 12310
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14292 11354 14320 11698
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 9518 14412 11086
rect 14476 10674 14504 12718
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 12442 14964 12650
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 15028 12306 15056 14486
rect 15120 13870 15148 16594
rect 15198 16280 15254 16289
rect 15198 16215 15200 16224
rect 15252 16215 15254 16224
rect 15200 16186 15252 16192
rect 15304 15688 15332 18663
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15212 15660 15332 15688
rect 15212 14793 15240 15660
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15304 15094 15332 15506
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15198 14784 15254 14793
rect 15198 14719 15254 14728
rect 15304 14482 15332 14894
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15120 13530 15148 13670
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15212 13462 15240 14214
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15304 12782 15332 13670
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14618 11996 14914 12016
rect 14674 11994 14698 11996
rect 14754 11994 14778 11996
rect 14834 11994 14858 11996
rect 14696 11942 14698 11994
rect 14760 11942 14772 11994
rect 14834 11942 14836 11994
rect 14674 11940 14698 11942
rect 14754 11940 14778 11942
rect 14834 11940 14858 11942
rect 14618 11920 14914 11940
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14752 11218 14780 11766
rect 15396 11354 15424 18566
rect 15488 18222 15516 19207
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16794 15516 17002
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15580 14929 15608 20726
rect 15566 14920 15622 14929
rect 15566 14855 15622 14864
rect 15672 14804 15700 23122
rect 15764 20466 15792 29242
rect 15856 29034 15884 29446
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 16040 28762 16068 28902
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 16132 28626 16160 30924
rect 16304 29096 16356 29102
rect 16304 29038 16356 29044
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 16120 28620 16172 28626
rect 16120 28562 16172 28568
rect 16040 27674 16068 28562
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15856 23526 15884 27474
rect 16028 26988 16080 26994
rect 16028 26930 16080 26936
rect 16040 25838 16068 26930
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 16028 25696 16080 25702
rect 16132 25684 16160 27814
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16224 25838 16252 26930
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 16132 25656 16252 25684
rect 16028 25638 16080 25644
rect 15934 24848 15990 24857
rect 15934 24783 15990 24792
rect 15948 24410 15976 24783
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 16040 23168 16068 25638
rect 16120 25152 16172 25158
rect 16120 25094 16172 25100
rect 16132 24274 16160 25094
rect 16224 24750 16252 25656
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16224 24070 16252 24686
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16212 23792 16264 23798
rect 16212 23734 16264 23740
rect 16224 23186 16252 23734
rect 15948 23140 16068 23168
rect 16212 23180 16264 23186
rect 15948 22166 15976 23140
rect 16212 23122 16264 23128
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15856 20806 15884 22034
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 15948 21078 15976 21354
rect 15936 21072 15988 21078
rect 15936 21014 15988 21020
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15764 19446 15792 20402
rect 15948 20398 15976 21014
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15764 19310 15792 19382
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15948 18834 15976 20334
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15764 17542 15792 17682
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15764 16658 15792 16934
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15948 16182 15976 18294
rect 16040 18086 16068 22986
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 16132 21622 16160 22442
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16026 16960 16082 16969
rect 16026 16895 16082 16904
rect 15936 16176 15988 16182
rect 15934 16144 15936 16153
rect 15988 16144 15990 16153
rect 15934 16079 15990 16088
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15764 14890 15792 15370
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15488 14776 15700 14804
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 14618 10908 14914 10928
rect 14674 10906 14698 10908
rect 14754 10906 14778 10908
rect 14834 10906 14858 10908
rect 14696 10854 14698 10906
rect 14760 10854 14772 10906
rect 14834 10854 14836 10906
rect 14674 10852 14698 10854
rect 14754 10852 14778 10854
rect 14834 10852 14858 10854
rect 14618 10832 14914 10852
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14618 9820 14914 9840
rect 14674 9818 14698 9820
rect 14754 9818 14778 9820
rect 14834 9818 14858 9820
rect 14696 9766 14698 9818
rect 14760 9766 14772 9818
rect 14834 9766 14836 9818
rect 14674 9764 14698 9766
rect 14754 9764 14778 9766
rect 14834 9764 14858 9766
rect 14618 9744 14914 9764
rect 15120 9602 15148 11018
rect 15212 10538 15240 11222
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 10606 15332 10950
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15396 10470 15424 11154
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 14936 9574 15148 9602
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14936 9042 14964 9574
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 9110 15056 9386
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14618 8732 14914 8752
rect 14674 8730 14698 8732
rect 14754 8730 14778 8732
rect 14834 8730 14858 8732
rect 14696 8678 14698 8730
rect 14760 8678 14772 8730
rect 14834 8678 14836 8730
rect 14674 8676 14698 8678
rect 14754 8676 14778 8678
rect 14834 8676 14858 8678
rect 14618 8656 14914 8676
rect 14186 8528 14242 8537
rect 14186 8463 14242 8472
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14200 6254 14228 8298
rect 14384 7954 14412 8366
rect 15304 8022 15332 8774
rect 15488 8090 15516 14776
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 12986 15608 13738
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15580 8430 15608 11290
rect 15672 9110 15700 14418
rect 15948 13530 15976 14486
rect 16040 13938 16068 16895
rect 16132 14482 16160 21286
rect 16224 19922 16252 21966
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16028 13932 16080 13938
rect 16224 13920 16252 17206
rect 16316 17066 16344 29038
rect 16396 28756 16448 28762
rect 16396 28698 16448 28704
rect 16408 27606 16436 28698
rect 16396 27600 16448 27606
rect 16396 27542 16448 27548
rect 16408 27062 16436 27542
rect 16592 27538 16620 30924
rect 17052 29102 17080 30924
rect 17972 29306 18000 30924
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17684 29096 17736 29102
rect 18052 29096 18104 29102
rect 17684 29038 17736 29044
rect 17972 29044 18052 29050
rect 17972 29038 18104 29044
rect 17592 28688 17644 28694
rect 17592 28630 17644 28636
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17236 28014 17264 28494
rect 17408 28484 17460 28490
rect 17408 28426 17460 28432
rect 17224 28008 17276 28014
rect 17224 27950 17276 27956
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 16948 27328 17000 27334
rect 16948 27270 17000 27276
rect 16396 27056 16448 27062
rect 16396 26998 16448 27004
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 16408 25974 16436 26862
rect 16672 26852 16724 26858
rect 16672 26794 16724 26800
rect 16580 26784 16632 26790
rect 16580 26726 16632 26732
rect 16396 25968 16448 25974
rect 16396 25910 16448 25916
rect 16408 22710 16436 25910
rect 16592 23186 16620 26726
rect 16684 26586 16712 26794
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 25362 16712 26522
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16408 19334 16436 21558
rect 16408 19306 16528 19334
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16316 15473 16344 15982
rect 16302 15464 16358 15473
rect 16302 15399 16358 15408
rect 16316 14550 16344 15399
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16028 13874 16080 13880
rect 16132 13892 16252 13920
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15750 12880 15806 12889
rect 15750 12815 15806 12824
rect 15764 12306 15792 12815
rect 15948 12617 15976 13126
rect 15934 12608 15990 12617
rect 15934 12543 15990 12552
rect 15842 12472 15898 12481
rect 15842 12407 15898 12416
rect 15856 12374 15884 12407
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15856 11898 15884 12106
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15948 11694 15976 12543
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16040 11082 16068 12242
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16132 10810 16160 13892
rect 16210 13832 16266 13841
rect 16210 13767 16266 13776
rect 16224 12442 16252 13767
rect 16316 13462 16344 14486
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16224 10742 16252 12378
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 8634 15792 8910
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14618 7644 14914 7664
rect 14674 7642 14698 7644
rect 14754 7642 14778 7644
rect 14834 7642 14858 7644
rect 14696 7590 14698 7642
rect 14760 7590 14772 7642
rect 14834 7590 14836 7642
rect 14674 7588 14698 7590
rect 14754 7588 14778 7590
rect 14834 7588 14858 7590
rect 14618 7568 14914 7588
rect 14618 6556 14914 6576
rect 14674 6554 14698 6556
rect 14754 6554 14778 6556
rect 14834 6554 14858 6556
rect 14696 6502 14698 6554
rect 14760 6502 14772 6554
rect 14834 6502 14836 6554
rect 14674 6500 14698 6502
rect 14754 6500 14778 6502
rect 14834 6500 14858 6502
rect 14618 6480 14914 6500
rect 14004 6248 14056 6254
rect 14002 6216 14004 6225
rect 14188 6248 14240 6254
rect 14056 6216 14058 6225
rect 14188 6190 14240 6196
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 14002 6151 14058 6160
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14016 4146 14044 5714
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14108 4486 14136 5170
rect 14384 4486 14412 6190
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5302 14504 6054
rect 14660 5642 14688 6122
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14618 5468 14914 5488
rect 14674 5466 14698 5468
rect 14754 5466 14778 5468
rect 14834 5466 14858 5468
rect 14696 5414 14698 5466
rect 14760 5414 14772 5466
rect 14834 5414 14836 5466
rect 14674 5412 14698 5414
rect 14754 5412 14778 5414
rect 14834 5412 14858 5414
rect 14618 5392 14914 5412
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4554 14504 4966
rect 15028 4758 15056 6054
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15120 5030 15148 5782
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 13924 3670 13952 4014
rect 14108 3942 14136 4014
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14384 3670 14412 4422
rect 14618 4380 14914 4400
rect 14674 4378 14698 4380
rect 14754 4378 14778 4380
rect 14834 4378 14858 4380
rect 14696 4326 14698 4378
rect 14760 4326 14772 4378
rect 14834 4326 14836 4378
rect 14674 4324 14698 4326
rect 14754 4324 14778 4326
rect 14834 4324 14858 4326
rect 14618 4304 14914 4324
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3194 13768 3334
rect 13924 3194 13952 3606
rect 14618 3292 14914 3312
rect 14674 3290 14698 3292
rect 14754 3290 14778 3292
rect 14834 3290 14858 3292
rect 14696 3238 14698 3290
rect 14760 3238 14772 3290
rect 14834 3238 14836 3290
rect 14674 3236 14698 3238
rect 14754 3236 14778 3238
rect 14834 3236 14858 3238
rect 14618 3216 14914 3236
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 15120 2990 15148 3946
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 13832 800 13860 2450
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13924 1902 13952 2246
rect 13912 1896 13964 1902
rect 13912 1838 13964 1844
rect 14292 800 14320 2450
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14618 2204 14914 2224
rect 14674 2202 14698 2204
rect 14754 2202 14778 2204
rect 14834 2202 14858 2204
rect 14696 2150 14698 2202
rect 14760 2150 14772 2202
rect 14834 2150 14836 2202
rect 14674 2148 14698 2150
rect 14754 2148 14778 2150
rect 14834 2148 14858 2150
rect 14618 2128 14914 2148
rect 15028 1834 15056 2314
rect 15016 1828 15068 1834
rect 15016 1770 15068 1776
rect 15212 800 15240 6190
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15304 4690 15332 5646
rect 15856 5166 15884 6190
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15304 4214 15332 4626
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15304 3534 15332 4150
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15474 3496 15530 3505
rect 15474 3431 15476 3440
rect 15528 3431 15530 3440
rect 15476 3402 15528 3408
rect 15672 800 15700 3538
rect 15948 2990 15976 6054
rect 16132 4049 16160 10406
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 7750 16344 8978
rect 16408 7818 16436 18022
rect 16500 17814 16528 19306
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16794 16528 16934
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16500 15638 16528 16730
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16500 12850 16528 13738
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16500 11286 16528 12786
rect 16592 12306 16620 18566
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16670 17640 16726 17649
rect 16670 17575 16672 17584
rect 16724 17575 16726 17584
rect 16672 17546 16724 17552
rect 16776 14550 16804 18090
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16684 12646 16712 13126
rect 16776 12730 16804 14486
rect 16868 14482 16896 14758
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16776 12702 16896 12730
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16592 11830 16620 12038
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16592 9042 16620 11562
rect 16776 11218 16804 12582
rect 16868 12170 16896 12702
rect 16960 12374 16988 27270
rect 17236 26450 17264 27950
rect 17420 27606 17448 28426
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 17512 27402 17540 28358
rect 17500 27396 17552 27402
rect 17500 27338 17552 27344
rect 17512 26926 17540 27338
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 17236 25838 17264 26386
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 17040 25220 17092 25226
rect 17040 25162 17092 25168
rect 17052 22234 17080 25162
rect 17236 23594 17264 25774
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17224 23588 17276 23594
rect 17224 23530 17276 23536
rect 17236 23050 17264 23530
rect 17328 23322 17356 25298
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17420 24138 17448 24686
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 24342 17540 24550
rect 17500 24336 17552 24342
rect 17500 24278 17552 24284
rect 17408 24132 17460 24138
rect 17408 24074 17460 24080
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17604 22574 17632 28630
rect 17696 27946 17724 29038
rect 17972 29022 18092 29038
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17696 27470 17724 27882
rect 17972 27878 18000 29022
rect 18144 28960 18196 28966
rect 18144 28902 18196 28908
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 27538 18000 27814
rect 18064 27674 18092 28562
rect 18156 28014 18184 28902
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 17960 27532 18012 27538
rect 17960 27474 18012 27480
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17696 24138 17724 27406
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17880 26518 17908 26726
rect 17868 26512 17920 26518
rect 17868 26454 17920 26460
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17696 23866 17724 24074
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17972 23526 18000 27474
rect 18340 26926 18368 27542
rect 18432 27538 18460 30924
rect 18892 29238 18920 30924
rect 19812 29238 19840 30924
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 18880 29232 18932 29238
rect 18880 29174 18932 29180
rect 19800 29232 19852 29238
rect 19800 29174 19852 29180
rect 19708 29164 19760 29170
rect 19708 29106 19760 29112
rect 18788 29028 18840 29034
rect 18788 28970 18840 28976
rect 18800 28150 18828 28970
rect 19172 28860 19468 28880
rect 19228 28858 19252 28860
rect 19308 28858 19332 28860
rect 19388 28858 19412 28860
rect 19250 28806 19252 28858
rect 19314 28806 19326 28858
rect 19388 28806 19390 28858
rect 19228 28804 19252 28806
rect 19308 28804 19332 28806
rect 19388 28804 19412 28806
rect 19172 28784 19468 28804
rect 18880 28416 18932 28422
rect 18880 28358 18932 28364
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18708 27130 18736 27270
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18800 26926 18828 28086
rect 18892 27606 18920 28358
rect 19720 28014 19748 29106
rect 20088 28626 20116 29514
rect 20272 28694 20300 30924
rect 20732 29306 20760 30924
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 21180 29300 21232 29306
rect 21180 29242 21232 29248
rect 20996 28960 21048 28966
rect 20996 28902 21048 28908
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 21008 28626 21036 28902
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 19172 27772 19468 27792
rect 19228 27770 19252 27772
rect 19308 27770 19332 27772
rect 19388 27770 19412 27772
rect 19250 27718 19252 27770
rect 19314 27718 19326 27770
rect 19388 27718 19390 27770
rect 19228 27716 19252 27718
rect 19308 27716 19332 27718
rect 19388 27716 19412 27718
rect 19172 27696 19468 27716
rect 18880 27600 18932 27606
rect 18880 27542 18932 27548
rect 18328 26920 18380 26926
rect 18328 26862 18380 26868
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18248 26586 18276 26794
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18604 26784 18656 26790
rect 18604 26726 18656 26732
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 18156 24750 18184 25298
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18340 24750 18368 25094
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 17960 23520 18012 23526
rect 17960 23462 18012 23468
rect 18432 23322 18460 23530
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 17880 22642 17908 23122
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17684 22568 17736 22574
rect 17684 22510 17736 22516
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 17052 21622 17080 22170
rect 17328 21894 17356 22510
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17420 22030 17448 22442
rect 17604 22234 17632 22510
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 17052 21010 17080 21422
rect 17132 21072 17184 21078
rect 17184 21020 17264 21026
rect 17132 21014 17264 21020
rect 17040 21004 17092 21010
rect 17144 20998 17264 21014
rect 17040 20946 17092 20952
rect 17052 15570 17080 20946
rect 17236 20330 17264 20998
rect 17328 20942 17356 21830
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 18737 17172 19110
rect 17130 18728 17186 18737
rect 17130 18663 17186 18672
rect 17236 16538 17264 20266
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17328 19514 17356 19858
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17420 18086 17448 21966
rect 17604 21622 17632 22170
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17202 17448 18022
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17328 16726 17356 16934
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17236 16510 17356 16538
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17052 14090 17080 15506
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17236 14600 17264 15370
rect 17328 15026 17356 16510
rect 17420 15978 17448 16934
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17236 14572 17356 14600
rect 17222 14512 17278 14521
rect 17222 14447 17224 14456
rect 17276 14447 17278 14456
rect 17224 14418 17276 14424
rect 17052 14062 17172 14090
rect 17040 13864 17092 13870
rect 17144 13852 17172 14062
rect 17144 13824 17264 13852
rect 17040 13806 17092 13812
rect 17052 13394 17080 13806
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 17052 12186 17080 13330
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16960 12158 17080 12186
rect 16868 11937 16896 12106
rect 16854 11928 16910 11937
rect 16854 11863 16910 11872
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16224 5302 16252 5714
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16118 4040 16174 4049
rect 16118 3975 16174 3984
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16040 2514 16068 2790
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16132 800 16160 3878
rect 16316 3097 16344 7686
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16408 6458 16436 6802
rect 16500 6662 16528 7278
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16408 6066 16436 6190
rect 16500 6186 16528 6598
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16408 6038 16528 6066
rect 16500 5710 16528 6038
rect 16592 5914 16620 7890
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 5166 16528 5646
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16592 5098 16620 5850
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16684 4010 16712 11018
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16776 3890 16804 11018
rect 16868 8838 16896 11766
rect 16960 11694 16988 12158
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16960 9518 16988 10678
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16960 6866 16988 8978
rect 17052 7546 17080 12038
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11082 17172 11630
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17144 10198 17172 11018
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17236 9110 17264 13824
rect 17328 13326 17356 14572
rect 17420 14482 17448 15302
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17512 14278 17540 21558
rect 17696 21078 17724 22510
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 17880 22098 17908 22374
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 18064 21434 18092 22374
rect 17972 21406 18092 21434
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 19446 17632 19654
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17604 18834 17632 19382
rect 17788 18834 17816 20742
rect 17972 20210 18000 21406
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 20398 18092 21286
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17972 20182 18092 20210
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17880 18766 17908 19314
rect 17868 18760 17920 18766
rect 17590 18728 17646 18737
rect 17868 18702 17920 18708
rect 17590 18663 17646 18672
rect 17604 14958 17632 18663
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17776 17196 17828 17202
rect 17880 17184 17908 18702
rect 18064 18358 18092 20182
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17828 17156 17908 17184
rect 17776 17138 17828 17144
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17604 14657 17632 14894
rect 17590 14648 17646 14657
rect 17590 14583 17646 14592
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17696 14090 17724 17138
rect 17512 14062 17724 14090
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17328 12442 17356 12718
rect 17420 12646 17448 12786
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17314 11928 17370 11937
rect 17314 11863 17370 11872
rect 17328 10674 17356 11863
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17420 11354 17448 11562
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9654 17356 10066
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16960 6186 16988 6802
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16684 3862 16804 3890
rect 16302 3088 16358 3097
rect 16302 3023 16358 3032
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16408 2514 16436 2994
rect 16684 2961 16712 3862
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16670 2952 16726 2961
rect 16670 2887 16726 2896
rect 16776 2650 16804 3538
rect 16868 2990 16896 6054
rect 16960 5778 16988 6122
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16960 4758 16988 5714
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16960 3398 16988 4014
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16960 2582 16988 3334
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 17052 800 17080 3538
rect 17144 2378 17172 7822
rect 17236 5574 17264 8366
rect 17328 7546 17356 9454
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17420 6338 17448 10950
rect 17328 6322 17448 6338
rect 17316 6316 17448 6322
rect 17368 6310 17448 6316
rect 17316 6258 17368 6264
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17420 5846 17448 6190
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17420 5166 17448 5782
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17236 4457 17264 4490
rect 17222 4448 17278 4457
rect 17222 4383 17278 4392
rect 17236 3058 17264 4383
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17512 2774 17540 14062
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17696 12918 17724 13126
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17604 12374 17632 12718
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17604 11014 17632 12174
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17604 9926 17632 10678
rect 17696 10266 17724 12242
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 8906 17632 9862
rect 17696 9518 17724 10202
rect 17788 9586 17816 17138
rect 17960 16992 18012 16998
rect 18052 16992 18104 16998
rect 17960 16934 18012 16940
rect 18050 16960 18052 16969
rect 18104 16960 18106 16969
rect 17972 16794 18000 16934
rect 18050 16895 18106 16904
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 16182 17908 16594
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17880 15434 17908 15982
rect 17972 15570 18000 16730
rect 18064 15978 18092 16730
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17960 15020 18012 15026
rect 17880 14980 17960 15008
rect 17880 10742 17908 14980
rect 17960 14962 18012 14968
rect 17958 14648 18014 14657
rect 17958 14583 18014 14592
rect 17972 13977 18000 14583
rect 18064 14482 18092 15302
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17958 13968 18014 13977
rect 17958 13903 18014 13912
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17972 13530 18000 13738
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18064 13258 18092 14214
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18156 12186 18184 22986
rect 18248 22574 18276 23122
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18248 22137 18276 22510
rect 18234 22128 18290 22137
rect 18234 22063 18290 22072
rect 18340 21962 18368 22510
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18432 22234 18460 22442
rect 18420 22228 18472 22234
rect 18420 22170 18472 22176
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18248 21593 18276 21626
rect 18234 21584 18290 21593
rect 18234 21519 18290 21528
rect 18236 21480 18288 21486
rect 18234 21448 18236 21457
rect 18288 21448 18290 21457
rect 18234 21383 18290 21392
rect 18248 21010 18276 21383
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18248 18970 18276 20334
rect 18340 19990 18368 21898
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18432 20874 18460 21626
rect 18524 21010 18552 26726
rect 18616 21486 18644 26726
rect 19172 26684 19468 26704
rect 19228 26682 19252 26684
rect 19308 26682 19332 26684
rect 19388 26682 19412 26684
rect 19250 26630 19252 26682
rect 19314 26630 19326 26682
rect 19388 26630 19390 26682
rect 19228 26628 19252 26630
rect 19308 26628 19332 26630
rect 19388 26628 19412 26630
rect 19172 26608 19468 26628
rect 18788 26580 18840 26586
rect 18788 26522 18840 26528
rect 18800 25362 18828 26522
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18708 24954 18736 25230
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18892 24750 18920 25638
rect 19172 25596 19468 25616
rect 19228 25594 19252 25596
rect 19308 25594 19332 25596
rect 19388 25594 19412 25596
rect 19250 25542 19252 25594
rect 19314 25542 19326 25594
rect 19388 25542 19390 25594
rect 19228 25540 19252 25542
rect 19308 25540 19332 25542
rect 19388 25540 19412 25542
rect 19172 25520 19468 25540
rect 19064 24880 19116 24886
rect 19064 24822 19116 24828
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18972 24676 19024 24682
rect 18972 24618 19024 24624
rect 18786 23352 18842 23361
rect 18696 23316 18748 23322
rect 18786 23287 18842 23296
rect 18696 23258 18748 23264
rect 18708 23225 18736 23258
rect 18800 23254 18828 23287
rect 18788 23248 18840 23254
rect 18694 23216 18750 23225
rect 18788 23190 18840 23196
rect 18694 23151 18750 23160
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18696 23112 18748 23118
rect 18892 23066 18920 23122
rect 18696 23054 18748 23060
rect 18708 21978 18736 23054
rect 18800 23038 18920 23066
rect 18800 22438 18828 23038
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18708 21950 18828 21978
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18420 20868 18472 20874
rect 18420 20810 18472 20816
rect 18432 20602 18460 20810
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 18616 20466 18644 21286
rect 18708 21010 18736 21830
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18708 19990 18736 20334
rect 18800 20262 18828 21950
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18340 19310 18368 19926
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18248 17066 18276 18362
rect 18432 18154 18460 19858
rect 18800 19836 18828 20198
rect 18708 19808 18828 19836
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18616 18290 18644 18770
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18234 16280 18290 16289
rect 18234 16215 18290 16224
rect 18248 16182 18276 16215
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18340 14958 18368 15914
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14550 18368 14758
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18234 13968 18290 13977
rect 18234 13903 18290 13912
rect 18248 13394 18276 13903
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18248 12889 18276 13330
rect 18234 12880 18290 12889
rect 18234 12815 18290 12824
rect 18340 12782 18368 13738
rect 18432 13190 18460 18090
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18616 16250 18644 17682
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18524 14793 18552 15030
rect 18510 14784 18566 14793
rect 18510 14719 18566 14728
rect 18510 14512 18566 14521
rect 18510 14447 18512 14456
rect 18564 14447 18566 14456
rect 18512 14418 18564 14424
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18248 12442 18276 12718
rect 18340 12617 18368 12718
rect 18326 12608 18382 12617
rect 18326 12543 18382 12552
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18156 12158 18368 12186
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 11354 18000 11630
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18064 11234 18092 11562
rect 18156 11558 18184 12038
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 17972 11218 18092 11234
rect 17960 11212 18092 11218
rect 18012 11206 18092 11212
rect 18340 11200 18368 12158
rect 18432 11218 18460 13126
rect 17960 11154 18012 11160
rect 18248 11172 18368 11200
rect 18420 11212 18472 11218
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 10266 17908 10542
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 9058 17724 9318
rect 17776 9104 17828 9110
rect 17696 9052 17776 9058
rect 17696 9046 17828 9052
rect 17696 9030 17816 9046
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17604 7410 17632 8298
rect 17696 7954 17724 9030
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17788 8566 17816 8774
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17788 7750 17816 8502
rect 17880 7954 17908 8842
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 18064 7886 18092 8366
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 6934 17632 7346
rect 17972 7342 18000 7686
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18064 7206 18092 7822
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 5284 17632 6870
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17696 6361 17724 6394
rect 17682 6352 17738 6361
rect 17682 6287 17738 6296
rect 17880 6254 17908 6666
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17684 5296 17736 5302
rect 17604 5256 17684 5284
rect 17684 5238 17736 5244
rect 17696 4690 17724 5238
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17972 4706 18000 5170
rect 17788 4690 18000 4706
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17776 4684 18000 4690
rect 17828 4678 18000 4684
rect 17776 4626 17828 4632
rect 17696 4214 17724 4626
rect 17684 4208 17736 4214
rect 17684 4150 17736 4156
rect 17972 4078 18000 4678
rect 18064 4486 18092 6802
rect 18248 6202 18276 11172
rect 18420 11154 18472 11160
rect 18432 11098 18460 11154
rect 18340 11070 18460 11098
rect 18340 10112 18368 11070
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10606 18460 10950
rect 18524 10674 18552 14418
rect 18616 13326 18644 15982
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18708 12434 18736 19808
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18800 17882 18828 19246
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18800 16726 18828 17818
rect 18892 17746 18920 22918
rect 18984 22148 19012 24618
rect 19076 22216 19104 24822
rect 19172 24508 19468 24528
rect 19228 24506 19252 24508
rect 19308 24506 19332 24508
rect 19388 24506 19412 24508
rect 19250 24454 19252 24506
rect 19314 24454 19326 24506
rect 19388 24454 19390 24506
rect 19228 24452 19252 24454
rect 19308 24452 19332 24454
rect 19388 24452 19412 24454
rect 19172 24432 19468 24452
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19536 23866 19564 24210
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19172 23420 19468 23440
rect 19228 23418 19252 23420
rect 19308 23418 19332 23420
rect 19388 23418 19412 23420
rect 19250 23366 19252 23418
rect 19314 23366 19326 23418
rect 19388 23366 19390 23418
rect 19228 23364 19252 23366
rect 19308 23364 19332 23366
rect 19388 23364 19412 23366
rect 19172 23344 19468 23364
rect 19154 23080 19210 23089
rect 19536 23050 19564 23802
rect 19154 23015 19210 23024
rect 19524 23044 19576 23050
rect 19168 22506 19196 23015
rect 19524 22986 19576 22992
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 19172 22332 19468 22352
rect 19228 22330 19252 22332
rect 19308 22330 19332 22332
rect 19388 22330 19412 22332
rect 19250 22278 19252 22330
rect 19314 22278 19326 22330
rect 19388 22278 19390 22330
rect 19228 22276 19252 22278
rect 19308 22276 19332 22278
rect 19388 22276 19412 22278
rect 19172 22256 19468 22276
rect 19076 22188 19196 22216
rect 18984 22120 19104 22148
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18984 21622 19012 21898
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18984 20466 19012 21422
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18984 17542 19012 19858
rect 19076 18426 19104 22120
rect 19168 21486 19196 22188
rect 19248 22160 19300 22166
rect 19248 22102 19300 22108
rect 19260 21962 19288 22102
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19156 21480 19208 21486
rect 19260 21457 19288 21626
rect 19156 21422 19208 21428
rect 19246 21448 19302 21457
rect 19246 21383 19302 21392
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19172 21244 19468 21264
rect 19228 21242 19252 21244
rect 19308 21242 19332 21244
rect 19388 21242 19412 21244
rect 19250 21190 19252 21242
rect 19314 21190 19326 21242
rect 19388 21190 19390 21242
rect 19228 21188 19252 21190
rect 19308 21188 19332 21190
rect 19388 21188 19412 21190
rect 19172 21168 19468 21188
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 20398 19380 20810
rect 19536 20398 19564 21286
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19628 20602 19656 20878
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19172 20156 19468 20176
rect 19228 20154 19252 20156
rect 19308 20154 19332 20156
rect 19388 20154 19412 20156
rect 19250 20102 19252 20154
rect 19314 20102 19326 20154
rect 19388 20102 19390 20154
rect 19228 20100 19252 20102
rect 19308 20100 19332 20102
rect 19388 20100 19412 20102
rect 19172 20080 19468 20100
rect 19172 19068 19468 19088
rect 19228 19066 19252 19068
rect 19308 19066 19332 19068
rect 19388 19066 19412 19068
rect 19250 19014 19252 19066
rect 19314 19014 19326 19066
rect 19388 19014 19390 19066
rect 19228 19012 19252 19014
rect 19308 19012 19332 19014
rect 19388 19012 19412 19014
rect 19172 18992 19468 19012
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18984 16046 19012 17478
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18616 12406 18736 12434
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18420 10124 18472 10130
rect 18340 10084 18420 10112
rect 18420 10066 18472 10072
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8090 18552 8774
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18524 7954 18552 8026
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18524 7002 18552 7890
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18248 6174 18552 6202
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18156 4146 18184 5170
rect 18432 5166 18460 5646
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18248 4282 18276 5034
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18248 3670 18276 3946
rect 18340 3942 18368 4150
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18064 3194 18092 3538
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18248 2922 18276 3334
rect 18432 3058 18460 4082
rect 18524 3505 18552 6174
rect 18510 3496 18566 3505
rect 18510 3431 18566 3440
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17512 2746 17724 2774
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17512 800 17540 2450
rect 17696 2106 17724 2746
rect 17684 2100 17736 2106
rect 17684 2042 17736 2048
rect 17972 800 18000 2790
rect 18616 2774 18644 12406
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18708 10606 18736 12106
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 9518 18736 10406
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8430 18736 8774
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 7954 18736 8230
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 6746 18736 7890
rect 18800 6866 18828 14962
rect 18892 14890 18920 15302
rect 18970 15056 19026 15065
rect 18970 14991 19026 15000
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18984 14414 19012 14991
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18892 13870 18920 14350
rect 18880 13864 18932 13870
rect 19076 13818 19104 18362
rect 19172 17980 19468 18000
rect 19228 17978 19252 17980
rect 19308 17978 19332 17980
rect 19388 17978 19412 17980
rect 19250 17926 19252 17978
rect 19314 17926 19326 17978
rect 19388 17926 19390 17978
rect 19228 17924 19252 17926
rect 19308 17924 19332 17926
rect 19388 17924 19412 17926
rect 19172 17904 19468 17924
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19168 17270 19196 17478
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 19614 17232 19670 17241
rect 19614 17167 19616 17176
rect 19668 17167 19670 17176
rect 19616 17138 19668 17144
rect 19172 16892 19468 16912
rect 19228 16890 19252 16892
rect 19308 16890 19332 16892
rect 19388 16890 19412 16892
rect 19250 16838 19252 16890
rect 19314 16838 19326 16890
rect 19388 16838 19390 16890
rect 19228 16836 19252 16838
rect 19308 16836 19332 16838
rect 19388 16836 19412 16838
rect 19172 16816 19468 16836
rect 19720 16794 19748 27950
rect 20088 26738 20116 28562
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 27606 20852 27814
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 20352 27464 20404 27470
rect 20916 27418 20944 28494
rect 20352 27406 20404 27412
rect 19904 26710 20116 26738
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19812 22030 19840 22374
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19812 18766 19840 19790
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19812 16658 19840 18702
rect 19904 17218 19932 26710
rect 20364 26450 20392 27406
rect 20824 27390 20944 27418
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20088 22574 20116 23122
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19996 21010 20024 22442
rect 20088 21962 20116 22510
rect 20456 22098 20484 23122
rect 20640 23050 20668 23530
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20548 22166 20576 22578
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 20088 21146 20116 21898
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 20180 20516 20208 21898
rect 20272 21350 20300 22034
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20548 21486 20576 21830
rect 20640 21486 20668 22374
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 19996 20488 20208 20516
rect 19996 19417 20024 20488
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 19982 19408 20038 19417
rect 19982 19343 20038 19352
rect 19996 18358 20024 19343
rect 20088 18970 20116 20266
rect 20364 19786 20392 20266
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20364 19378 20392 19722
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19984 18216 20036 18222
rect 19982 18184 19984 18193
rect 20036 18184 20038 18193
rect 19982 18119 20038 18128
rect 20088 17882 20116 18770
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18222 20300 18566
rect 20364 18222 20392 19314
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20272 17746 20300 18158
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19904 17190 20208 17218
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19172 15804 19468 15824
rect 19228 15802 19252 15804
rect 19308 15802 19332 15804
rect 19388 15802 19412 15804
rect 19250 15750 19252 15802
rect 19314 15750 19326 15802
rect 19388 15750 19390 15802
rect 19228 15748 19252 15750
rect 19308 15748 19332 15750
rect 19388 15748 19412 15750
rect 19172 15728 19468 15748
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19172 14716 19468 14736
rect 19228 14714 19252 14716
rect 19308 14714 19332 14716
rect 19388 14714 19412 14716
rect 19250 14662 19252 14714
rect 19314 14662 19326 14714
rect 19388 14662 19390 14714
rect 19228 14660 19252 14662
rect 19308 14660 19332 14662
rect 19388 14660 19412 14662
rect 19172 14640 19468 14660
rect 18880 13806 18932 13812
rect 18984 13790 19104 13818
rect 18984 13530 19012 13790
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19076 13462 19104 13670
rect 19172 13628 19468 13648
rect 19228 13626 19252 13628
rect 19308 13626 19332 13628
rect 19388 13626 19412 13628
rect 19250 13574 19252 13626
rect 19314 13574 19326 13626
rect 19388 13574 19390 13626
rect 19228 13572 19252 13574
rect 19308 13572 19332 13574
rect 19388 13572 19412 13574
rect 19172 13552 19468 13572
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18892 12986 18920 13330
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18984 12481 19012 13194
rect 18970 12472 19026 12481
rect 18970 12407 19026 12416
rect 19076 12306 19104 13398
rect 19172 12540 19468 12560
rect 19228 12538 19252 12540
rect 19308 12538 19332 12540
rect 19388 12538 19412 12540
rect 19250 12486 19252 12538
rect 19314 12486 19326 12538
rect 19388 12486 19390 12538
rect 19228 12484 19252 12486
rect 19308 12484 19332 12486
rect 19388 12484 19412 12486
rect 19172 12464 19468 12484
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19172 11452 19468 11472
rect 19228 11450 19252 11452
rect 19308 11450 19332 11452
rect 19388 11450 19412 11452
rect 19250 11398 19252 11450
rect 19314 11398 19326 11450
rect 19388 11398 19390 11450
rect 19228 11396 19252 11398
rect 19308 11396 19332 11398
rect 19388 11396 19412 11398
rect 19172 11376 19468 11396
rect 19172 10364 19468 10384
rect 19228 10362 19252 10364
rect 19308 10362 19332 10364
rect 19388 10362 19412 10364
rect 19250 10310 19252 10362
rect 19314 10310 19326 10362
rect 19388 10310 19390 10362
rect 19228 10308 19252 10310
rect 19308 10308 19332 10310
rect 19388 10308 19412 10310
rect 19172 10288 19468 10308
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18708 6718 18828 6746
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18708 4622 18736 5102
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18708 4078 18736 4558
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18800 2774 18828 6718
rect 18892 3754 18920 10066
rect 19536 9654 19564 14894
rect 19628 14550 19656 15982
rect 19708 15972 19760 15978
rect 19708 15914 19760 15920
rect 19720 14929 19748 15914
rect 20088 15638 20116 16390
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 19890 15328 19946 15337
rect 19890 15263 19946 15272
rect 19904 14958 19932 15263
rect 20088 14958 20116 15574
rect 19892 14952 19944 14958
rect 19706 14920 19762 14929
rect 19892 14894 19944 14900
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19706 14855 19762 14864
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19628 12782 19656 14486
rect 19720 13938 19748 14758
rect 19996 14090 20024 14826
rect 19904 14062 20024 14090
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19720 12434 19748 12718
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19812 12442 19840 12650
rect 19628 12406 19748 12434
rect 19800 12436 19852 12442
rect 19628 12238 19656 12406
rect 19800 12378 19852 12384
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19628 11558 19656 12174
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19628 11082 19656 11494
rect 19812 11150 19840 12378
rect 19904 11286 19932 14062
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20088 12434 20116 13874
rect 19996 12406 20116 12434
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19628 10674 19656 11018
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 8634 19012 9454
rect 19172 9276 19468 9296
rect 19228 9274 19252 9276
rect 19308 9274 19332 9276
rect 19388 9274 19412 9276
rect 19250 9222 19252 9274
rect 19314 9222 19326 9274
rect 19388 9222 19390 9274
rect 19228 9220 19252 9222
rect 19308 9220 19332 9222
rect 19388 9220 19412 9222
rect 19172 9200 19468 9220
rect 19628 8838 19656 10610
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19720 8906 19748 9590
rect 19812 9042 19840 11086
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19904 9586 19932 9998
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19904 9110 19932 9386
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19892 8968 19944 8974
rect 19890 8936 19892 8945
rect 19944 8936 19946 8945
rect 19708 8900 19760 8906
rect 19890 8871 19946 8880
rect 19708 8842 19760 8848
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18970 8528 19026 8537
rect 18970 8463 19026 8472
rect 18984 8090 19012 8463
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18984 7478 19012 7890
rect 19076 7750 19104 8366
rect 19172 8188 19468 8208
rect 19228 8186 19252 8188
rect 19308 8186 19332 8188
rect 19388 8186 19412 8188
rect 19250 8134 19252 8186
rect 19314 8134 19326 8186
rect 19388 8134 19390 8186
rect 19228 8132 19252 8134
rect 19308 8132 19332 8134
rect 19388 8132 19412 8134
rect 19172 8112 19468 8132
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19720 7546 19748 8842
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 18972 7472 19024 7478
rect 19996 7426 20024 12406
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20088 8498 20116 11630
rect 20180 8634 20208 17190
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20272 16658 20300 17070
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20456 16046 20484 20946
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20640 19310 20668 20334
rect 20732 19514 20760 20946
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20732 19242 20760 19450
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20548 18426 20576 18770
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20548 15586 20576 18090
rect 20640 16250 20668 18158
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20732 17270 20760 17750
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20718 17096 20774 17105
rect 20718 17031 20774 17040
rect 20732 16998 20760 17031
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20456 15558 20576 15586
rect 20272 15094 20300 15506
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20272 12918 20300 13806
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20456 12730 20484 15558
rect 20640 14482 20668 16186
rect 20824 15910 20852 27390
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 20916 25498 20944 25774
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20902 22128 20958 22137
rect 20902 22063 20958 22072
rect 20916 21554 20944 22063
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 21008 21078 21036 28562
rect 21088 25764 21140 25770
rect 21088 25706 21140 25712
rect 21100 24682 21128 25706
rect 21088 24676 21140 24682
rect 21088 24618 21140 24624
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 20904 19304 20956 19310
rect 20956 19264 21036 19292
rect 20904 19246 20956 19252
rect 21008 18834 21036 19264
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 21008 18426 21036 18770
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21008 18193 21036 18362
rect 20994 18184 21050 18193
rect 20994 18119 21050 18128
rect 21100 17066 21128 24618
rect 21192 23322 21220 29242
rect 21284 28014 21312 29446
rect 21652 29102 21680 30924
rect 22112 29306 22140 30924
rect 22100 29300 22152 29306
rect 22100 29242 22152 29248
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 21732 28076 21784 28082
rect 21732 28018 21784 28024
rect 21272 28008 21324 28014
rect 21272 27950 21324 27956
rect 21640 28008 21692 28014
rect 21640 27950 21692 27956
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21652 26738 21680 27950
rect 21744 27402 21772 28018
rect 22572 28014 22600 30924
rect 23492 28626 23520 30924
rect 23952 29594 23980 30924
rect 23952 29566 24164 29594
rect 23726 29404 24022 29424
rect 23782 29402 23806 29404
rect 23862 29402 23886 29404
rect 23942 29402 23966 29404
rect 23804 29350 23806 29402
rect 23868 29350 23880 29402
rect 23942 29350 23944 29402
rect 23782 29348 23806 29350
rect 23862 29348 23886 29350
rect 23942 29348 23966 29350
rect 23726 29328 24022 29348
rect 23756 29028 23808 29034
rect 23756 28970 23808 28976
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23768 28558 23796 28970
rect 23756 28552 23808 28558
rect 23756 28494 23808 28500
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 21732 27396 21784 27402
rect 21732 27338 21784 27344
rect 21744 26926 21772 27338
rect 21732 26920 21784 26926
rect 21732 26862 21784 26868
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21468 26042 21496 26386
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21270 23624 21326 23633
rect 21270 23559 21326 23568
rect 21284 23526 21312 23559
rect 21468 23526 21496 24686
rect 21560 23594 21588 26726
rect 21652 26710 21772 26738
rect 21548 23588 21600 23594
rect 21548 23530 21600 23536
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21468 23118 21496 23462
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21376 22574 21404 22918
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 21284 20874 21312 22442
rect 21468 22166 21496 22510
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 21560 22098 21588 23054
rect 21652 22574 21680 23122
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19990 21220 20198
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21376 18086 21404 19178
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21546 17232 21602 17241
rect 21546 17167 21602 17176
rect 21560 17134 21588 17167
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16726 20944 16934
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 21100 16250 21128 17002
rect 21468 16794 21496 17070
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20810 15736 20866 15745
rect 20810 15671 20866 15680
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 14482 20760 15302
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20824 14414 20852 15671
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20272 12702 20484 12730
rect 20272 11762 20300 12702
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20364 11642 20392 12582
rect 20272 11614 20392 11642
rect 20272 9654 20300 11614
rect 20548 11506 20576 14282
rect 20916 13870 20944 15914
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20640 12646 20668 13806
rect 21008 13802 21036 15914
rect 21284 14958 21312 16186
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21362 14920 21418 14929
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20732 11830 20760 12242
rect 20720 11824 20772 11830
rect 20824 11801 20852 13194
rect 20720 11766 20772 11772
rect 20810 11792 20866 11801
rect 20810 11727 20866 11736
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20640 11506 20668 11630
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20364 11478 20668 11506
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20260 9512 20312 9518
rect 20364 9500 20392 11478
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20456 10266 20484 11154
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20312 9472 20392 9500
rect 20260 9454 20312 9460
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20180 8430 20208 8570
rect 20272 8566 20300 9454
rect 20456 9110 20484 10202
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20548 9178 20576 10066
rect 20640 9722 20668 11290
rect 20720 11212 20772 11218
rect 20824 11200 20852 11562
rect 20916 11218 20944 13670
rect 21100 13462 21128 14894
rect 21362 14855 21364 14864
rect 21416 14855 21418 14864
rect 21364 14826 21416 14832
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 21008 11354 21036 12650
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20772 11172 20852 11200
rect 20720 11154 20772 11160
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20732 9654 20760 10474
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20824 8650 20852 11172
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20916 11014 20944 11154
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20902 9616 20958 9625
rect 20902 9551 20958 9560
rect 20916 9518 20944 9551
rect 21008 9518 21036 10406
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 20732 8622 20852 8650
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 20088 7546 20116 7890
rect 20180 7886 20208 8366
rect 20732 8294 20760 8622
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 21100 8090 21128 13262
rect 21468 12434 21496 16730
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21652 14550 21680 15030
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21468 12406 21588 12434
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21192 11898 21220 12242
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21178 11792 21234 11801
rect 21178 11727 21234 11736
rect 21192 11694 21220 11727
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21284 11257 21312 12310
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21468 11286 21496 12242
rect 21560 11914 21588 12406
rect 21652 12306 21680 12582
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21560 11886 21680 11914
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21456 11280 21508 11286
rect 21270 11248 21326 11257
rect 21456 11222 21508 11228
rect 21270 11183 21326 11192
rect 21560 11082 21588 11698
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20902 7984 20958 7993
rect 21192 7954 21220 8230
rect 20902 7919 20904 7928
rect 20956 7919 20958 7928
rect 21180 7948 21232 7954
rect 20904 7890 20956 7896
rect 21180 7890 21232 7896
rect 20168 7880 20220 7886
rect 21272 7880 21324 7886
rect 20168 7822 20220 7828
rect 20258 7848 20314 7857
rect 21272 7822 21324 7828
rect 20258 7783 20314 7792
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 18972 7414 19024 7420
rect 19904 7398 20024 7426
rect 19172 7100 19468 7120
rect 19228 7098 19252 7100
rect 19308 7098 19332 7100
rect 19388 7098 19412 7100
rect 19250 7046 19252 7098
rect 19314 7046 19326 7098
rect 19388 7046 19390 7098
rect 19228 7044 19252 7046
rect 19308 7044 19332 7046
rect 19388 7044 19412 7046
rect 19172 7024 19468 7044
rect 19172 6012 19468 6032
rect 19228 6010 19252 6012
rect 19308 6010 19332 6012
rect 19388 6010 19412 6012
rect 19250 5958 19252 6010
rect 19314 5958 19326 6010
rect 19388 5958 19390 6010
rect 19228 5956 19252 5958
rect 19308 5956 19332 5958
rect 19388 5956 19412 5958
rect 19172 5936 19468 5956
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19524 5092 19576 5098
rect 19524 5034 19576 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18984 4214 19012 4490
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 19076 4078 19104 4966
rect 19172 4924 19468 4944
rect 19228 4922 19252 4924
rect 19308 4922 19332 4924
rect 19388 4922 19412 4924
rect 19250 4870 19252 4922
rect 19314 4870 19326 4922
rect 19388 4870 19390 4922
rect 19228 4868 19252 4870
rect 19308 4868 19332 4870
rect 19388 4868 19412 4870
rect 19172 4848 19468 4868
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19536 3942 19564 5034
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19172 3836 19468 3856
rect 19228 3834 19252 3836
rect 19308 3834 19332 3836
rect 19388 3834 19412 3836
rect 19250 3782 19252 3834
rect 19314 3782 19326 3834
rect 19388 3782 19390 3834
rect 19228 3780 19252 3782
rect 19308 3780 19332 3782
rect 19388 3780 19412 3782
rect 19172 3760 19468 3780
rect 18892 3726 19012 3754
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18432 2746 18644 2774
rect 18708 2746 18828 2774
rect 18432 2582 18460 2746
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18708 1766 18736 2746
rect 18696 1760 18748 1766
rect 18696 1702 18748 1708
rect 18892 800 18920 3538
rect 18984 3398 19012 3726
rect 19154 3632 19210 3641
rect 19154 3567 19210 3576
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 19168 3194 19196 3567
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19331 3052 19383 3058
rect 19331 2994 19383 3000
rect 19352 2961 19380 2994
rect 19338 2952 19394 2961
rect 19338 2887 19394 2896
rect 19172 2748 19468 2768
rect 19228 2746 19252 2748
rect 19308 2746 19332 2748
rect 19388 2746 19412 2748
rect 19250 2694 19252 2746
rect 19314 2694 19326 2746
rect 19388 2694 19390 2746
rect 19228 2692 19252 2694
rect 19308 2692 19332 2694
rect 19388 2692 19412 2694
rect 19172 2672 19468 2692
rect 19628 2582 19656 5510
rect 19708 4752 19760 4758
rect 19706 4720 19708 4729
rect 19760 4720 19762 4729
rect 19706 4655 19762 4664
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 19720 1442 19748 3674
rect 19352 1414 19748 1442
rect 19352 800 19380 1414
rect 19812 800 19840 5714
rect 19904 2990 19932 7398
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19996 5030 20024 7278
rect 20272 6934 20300 7783
rect 21180 7404 21232 7410
rect 21284 7392 21312 7822
rect 21232 7364 21312 7392
rect 21180 7346 21232 7352
rect 20536 7336 20588 7342
rect 21456 7336 21508 7342
rect 20536 7278 20588 7284
rect 21284 7296 21456 7324
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20548 6254 20576 7278
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6254 20852 6598
rect 21100 6458 21128 6802
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21284 6254 21312 7296
rect 21456 7278 21508 7284
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 20548 5846 20576 6190
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20456 5030 20484 5714
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 19996 4214 20024 4966
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 20180 3942 20208 4626
rect 20272 4486 20300 4694
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20258 3768 20314 3777
rect 20258 3703 20314 3712
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19996 2650 20024 3538
rect 20272 3534 20300 3703
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20074 3088 20130 3097
rect 20074 3023 20130 3032
rect 20088 2990 20116 3023
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19996 2446 20024 2586
rect 20180 2582 20208 2858
rect 20364 2854 20392 4422
rect 20456 3670 20484 4966
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20548 3602 20576 5782
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21008 4826 21036 5102
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20640 4729 20668 4762
rect 20626 4720 20682 4729
rect 20626 4655 20682 4664
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 20718 4176 20774 4185
rect 20718 4111 20720 4120
rect 20772 4111 20774 4120
rect 20720 4082 20772 4088
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 20456 2961 20484 3402
rect 20442 2952 20498 2961
rect 20442 2887 20498 2896
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20168 2576 20220 2582
rect 20168 2518 20220 2524
rect 20456 2514 20484 2887
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20548 2378 20576 3538
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 2650 20668 2790
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 20732 800 20760 2926
rect 21100 1442 21128 4014
rect 21192 3738 21220 4626
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 21284 3602 21312 6190
rect 21560 5302 21588 9318
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21652 4146 21680 11886
rect 21744 8430 21772 26710
rect 21836 25226 21864 26862
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22296 25838 22324 26522
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22192 25356 22244 25362
rect 22192 25298 22244 25304
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 22100 24880 22152 24886
rect 22100 24822 22152 24828
rect 22112 24274 22140 24822
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 22204 24154 22232 25298
rect 22112 24138 22232 24154
rect 22100 24132 22232 24138
rect 22152 24126 22232 24132
rect 22100 24074 22152 24080
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22204 22710 22232 24006
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21928 22166 21956 22578
rect 21916 22160 21968 22166
rect 21916 22102 21968 22108
rect 22296 22094 22324 25638
rect 22204 22066 22324 22094
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21836 20330 21864 20946
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21836 20058 21864 20266
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 22204 17542 22232 22066
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22204 17202 22232 17478
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21928 15638 21956 15914
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 21916 15360 21968 15366
rect 22112 15337 22140 15370
rect 21916 15302 21968 15308
rect 22098 15328 22154 15337
rect 21824 14476 21876 14482
rect 21928 14464 21956 15302
rect 22098 15263 22154 15272
rect 22112 15094 22140 15263
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22204 14929 22232 17138
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22190 14920 22246 14929
rect 22190 14855 22246 14864
rect 22296 14618 22324 15846
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 21876 14436 21956 14464
rect 21824 14418 21876 14424
rect 21928 12850 21956 14436
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 22112 12442 22140 13330
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22006 11792 22062 11801
rect 22006 11727 22062 11736
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21836 8906 21864 8978
rect 21928 8974 21956 10950
rect 22020 9625 22048 11727
rect 22112 11626 22140 12378
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22006 9616 22062 9625
rect 22006 9551 22062 9560
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 22020 8838 22048 9551
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22112 8616 22140 9046
rect 21928 8588 22140 8616
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21836 7410 21864 7958
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21192 2582 21220 3334
rect 21284 2650 21312 3538
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21180 2576 21232 2582
rect 21180 2518 21232 2524
rect 21100 1414 21220 1442
rect 21192 800 21220 1414
rect 21652 800 21680 2790
rect 21928 1834 21956 8588
rect 22204 8362 22232 11222
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22112 7274 22140 7890
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5098 22140 6054
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22020 3670 22048 4014
rect 22008 3664 22060 3670
rect 22008 3606 22060 3612
rect 22020 2650 22048 3606
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22204 1902 22232 8298
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22296 5030 22324 5306
rect 22388 5098 22416 27814
rect 22664 24562 22692 28358
rect 23726 28316 24022 28336
rect 23782 28314 23806 28316
rect 23862 28314 23886 28316
rect 23942 28314 23966 28316
rect 23804 28262 23806 28314
rect 23868 28262 23880 28314
rect 23942 28262 23944 28314
rect 23782 28260 23806 28262
rect 23862 28260 23886 28262
rect 23942 28260 23966 28262
rect 23726 28240 24022 28260
rect 24136 28014 24164 29566
rect 24412 28694 24440 30924
rect 24584 28960 24636 28966
rect 24584 28902 24636 28908
rect 24400 28688 24452 28694
rect 24400 28630 24452 28636
rect 24216 28620 24268 28626
rect 24216 28562 24268 28568
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 23726 27228 24022 27248
rect 23782 27226 23806 27228
rect 23862 27226 23886 27228
rect 23942 27226 23966 27228
rect 23804 27174 23806 27226
rect 23868 27174 23880 27226
rect 23942 27174 23944 27226
rect 23782 27172 23806 27174
rect 23862 27172 23886 27174
rect 23942 27172 23966 27174
rect 23726 27152 24022 27172
rect 22928 26920 22980 26926
rect 22928 26862 22980 26868
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 22848 25838 22876 26318
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 22940 25702 22968 26862
rect 23296 26852 23348 26858
rect 23296 26794 23348 26800
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 22928 25696 22980 25702
rect 22928 25638 22980 25644
rect 23216 24750 23244 26726
rect 23308 26586 23336 26794
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 23400 26518 23428 26726
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23726 26140 24022 26160
rect 23782 26138 23806 26140
rect 23862 26138 23886 26140
rect 23942 26138 23966 26140
rect 23804 26086 23806 26138
rect 23868 26086 23880 26138
rect 23942 26086 23944 26138
rect 23782 26084 23806 26086
rect 23862 26084 23886 26086
rect 23942 26084 23966 26086
rect 23726 26064 24022 26084
rect 24228 26042 24256 28562
rect 24596 28014 24624 28902
rect 25044 28620 25096 28626
rect 25044 28562 25096 28568
rect 24584 28008 24636 28014
rect 24412 27968 24584 27996
rect 24308 27532 24360 27538
rect 24308 27474 24360 27480
rect 24320 26926 24348 27474
rect 24308 26920 24360 26926
rect 24308 26862 24360 26868
rect 24320 26586 24348 26862
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24216 26036 24268 26042
rect 24216 25978 24268 25984
rect 23388 25764 23440 25770
rect 23388 25706 23440 25712
rect 23400 25498 23428 25706
rect 24124 25696 24176 25702
rect 24124 25638 24176 25644
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23296 25424 23348 25430
rect 23296 25366 23348 25372
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23308 24682 23336 25366
rect 23726 25052 24022 25072
rect 23782 25050 23806 25052
rect 23862 25050 23886 25052
rect 23942 25050 23966 25052
rect 23804 24998 23806 25050
rect 23868 24998 23880 25050
rect 23942 24998 23944 25050
rect 23782 24996 23806 24998
rect 23862 24996 23886 24998
rect 23942 24996 23966 24998
rect 23726 24976 24022 24996
rect 24136 24750 24164 25638
rect 24228 25362 24256 25978
rect 24216 25356 24268 25362
rect 24216 25298 24268 25304
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 23296 24676 23348 24682
rect 23296 24618 23348 24624
rect 22572 24534 22692 24562
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22480 21146 22508 24210
rect 22572 22522 22600 24534
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22664 23730 22692 24346
rect 22940 24274 22968 24550
rect 22928 24268 22980 24274
rect 22928 24210 22980 24216
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 23032 23746 23060 24006
rect 23204 23792 23256 23798
rect 23032 23740 23204 23746
rect 23032 23734 23256 23740
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 23032 23718 23244 23734
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22756 23322 22784 23598
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 22572 22506 22692 22522
rect 22572 22500 22704 22506
rect 22572 22494 22652 22500
rect 22652 22442 22704 22448
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22572 21894 22600 22374
rect 22664 22234 22692 22442
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22572 21010 22600 21830
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22664 21146 22692 21422
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22480 19174 22508 20810
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 22664 19446 22692 19994
rect 22940 19990 22968 22170
rect 23032 21690 23060 23718
rect 23308 22794 23336 24618
rect 23400 24614 23428 24686
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23726 23964 24022 23984
rect 23782 23962 23806 23964
rect 23862 23962 23886 23964
rect 23942 23962 23966 23964
rect 23804 23910 23806 23962
rect 23868 23910 23880 23962
rect 23942 23910 23944 23962
rect 23782 23908 23806 23910
rect 23862 23908 23886 23910
rect 23942 23908 23966 23910
rect 23726 23888 24022 23908
rect 23940 23656 23992 23662
rect 24136 23644 24164 24686
rect 23992 23616 24164 23644
rect 23940 23598 23992 23604
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23216 22766 23336 22794
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 23124 22166 23152 22374
rect 23112 22160 23164 22166
rect 23112 22102 23164 22108
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 23032 21078 23060 21626
rect 23216 21622 23244 22766
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23020 21072 23072 21078
rect 23020 21014 23072 21020
rect 23124 20398 23152 21286
rect 23308 20398 23336 22646
rect 23492 22642 23520 22986
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23492 22098 23520 22578
rect 23584 22098 23612 23462
rect 23952 23050 23980 23598
rect 24216 23588 24268 23594
rect 24216 23530 24268 23536
rect 24124 23180 24176 23186
rect 24124 23122 24176 23128
rect 23940 23044 23992 23050
rect 23940 22986 23992 22992
rect 23726 22876 24022 22896
rect 23782 22874 23806 22876
rect 23862 22874 23886 22876
rect 23942 22874 23966 22876
rect 23804 22822 23806 22874
rect 23868 22822 23880 22874
rect 23942 22822 23944 22874
rect 23782 22820 23806 22822
rect 23862 22820 23886 22822
rect 23942 22820 23966 22822
rect 23726 22800 24022 22820
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 22098 23980 22646
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 23860 21962 23888 22034
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23112 20392 23164 20398
rect 23112 20334 23164 20340
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23400 20330 23428 21898
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23584 21486 23612 21830
rect 23726 21788 24022 21808
rect 23782 21786 23806 21788
rect 23862 21786 23886 21788
rect 23942 21786 23966 21788
rect 23804 21734 23806 21786
rect 23868 21734 23880 21786
rect 23942 21734 23944 21786
rect 23782 21732 23806 21734
rect 23862 21732 23886 21734
rect 23942 21732 23966 21734
rect 23726 21712 24022 21732
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23480 20800 23532 20806
rect 23676 20788 23704 21558
rect 23952 21486 23980 21558
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 24136 20890 24164 23122
rect 24228 21690 24256 23530
rect 24308 23248 24360 23254
rect 24308 23190 24360 23196
rect 24320 22982 24348 23190
rect 24308 22976 24360 22982
rect 24308 22918 24360 22924
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24320 21486 24348 22918
rect 24412 22234 24440 27968
rect 24584 27950 24636 27956
rect 24676 27872 24728 27878
rect 24676 27814 24728 27820
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24308 21480 24360 21486
rect 24308 21422 24360 21428
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 24228 20992 24256 21354
rect 24412 21146 24440 22170
rect 24596 21554 24624 22510
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24228 20964 24440 20992
rect 24136 20862 24348 20890
rect 23480 20742 23532 20748
rect 23584 20760 23704 20788
rect 24124 20800 24176 20806
rect 23492 20466 23520 20742
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23584 19990 23612 20760
rect 24124 20742 24176 20748
rect 23726 20700 24022 20720
rect 23782 20698 23806 20700
rect 23862 20698 23886 20700
rect 23942 20698 23966 20700
rect 23804 20646 23806 20698
rect 23868 20646 23880 20698
rect 23942 20646 23944 20698
rect 23782 20644 23806 20646
rect 23862 20644 23886 20646
rect 23942 20644 23966 20646
rect 23726 20624 24022 20644
rect 24136 20398 24164 20742
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22572 18086 22600 19178
rect 22756 18834 22784 19858
rect 23216 19514 23244 19858
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 22928 19168 22980 19174
rect 22928 19110 22980 19116
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22940 18834 22968 19110
rect 23032 18902 23060 19110
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 23216 18834 23244 19450
rect 23296 19236 23348 19242
rect 23296 19178 23348 19184
rect 23308 18970 23336 19178
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 22940 18578 22968 18770
rect 22940 18550 23060 18578
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22480 16658 22508 16934
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22572 16590 22600 18022
rect 22742 17096 22798 17105
rect 22742 17031 22744 17040
rect 22796 17031 22798 17040
rect 22744 17002 22796 17008
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22480 14618 22508 14758
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22572 12442 22600 13262
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22664 11218 22692 12174
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22756 8634 22784 11018
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22940 10962 22968 14894
rect 23032 11082 23060 18550
rect 23492 17814 23520 19858
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23584 19242 23612 19654
rect 23726 19612 24022 19632
rect 23782 19610 23806 19612
rect 23862 19610 23886 19612
rect 23942 19610 23966 19612
rect 23804 19558 23806 19610
rect 23868 19558 23880 19610
rect 23942 19558 23944 19610
rect 23782 19556 23806 19558
rect 23862 19556 23886 19558
rect 23942 19556 23966 19558
rect 23726 19536 24022 19556
rect 23572 19236 23624 19242
rect 23572 19178 23624 19184
rect 24136 18698 24164 19926
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 23726 18524 24022 18544
rect 23782 18522 23806 18524
rect 23862 18522 23886 18524
rect 23942 18522 23966 18524
rect 23804 18470 23806 18522
rect 23868 18470 23880 18522
rect 23942 18470 23944 18522
rect 23782 18468 23806 18470
rect 23862 18468 23886 18470
rect 23942 18468 23966 18470
rect 23726 18448 24022 18468
rect 24320 18222 24348 20862
rect 24412 18986 24440 20964
rect 24504 19174 24532 21422
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24596 19854 24624 20946
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24596 19174 24624 19790
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24412 18958 24532 18986
rect 24400 18828 24452 18834
rect 24400 18770 24452 18776
rect 24412 18426 24440 18770
rect 24504 18766 24532 18958
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24308 18216 24360 18222
rect 24308 18158 24360 18164
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23124 16726 23152 16934
rect 23112 16720 23164 16726
rect 23112 16662 23164 16668
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23400 15722 23428 16118
rect 23492 16046 23520 17750
rect 23726 17436 24022 17456
rect 23782 17434 23806 17436
rect 23862 17434 23886 17436
rect 23942 17434 23966 17436
rect 23804 17382 23806 17434
rect 23868 17382 23880 17434
rect 23942 17382 23944 17434
rect 23782 17380 23806 17382
rect 23862 17380 23886 17382
rect 23942 17380 23966 17382
rect 23726 17360 24022 17380
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23952 16794 23980 17070
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 24492 16788 24544 16794
rect 24492 16730 24544 16736
rect 23726 16348 24022 16368
rect 23782 16346 23806 16348
rect 23862 16346 23886 16348
rect 23942 16346 23966 16348
rect 23804 16294 23806 16346
rect 23868 16294 23880 16346
rect 23942 16294 23944 16346
rect 23782 16292 23806 16294
rect 23862 16292 23886 16294
rect 23942 16292 23966 16294
rect 23726 16272 24022 16292
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23308 15706 23428 15722
rect 23308 15700 23440 15706
rect 23308 15694 23388 15700
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23216 14482 23244 15098
rect 23308 14958 23336 15694
rect 23388 15642 23440 15648
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23400 15162 23428 15506
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23480 15088 23532 15094
rect 23400 15036 23480 15042
rect 23400 15030 23532 15036
rect 23400 15014 23520 15030
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 23124 14074 23152 14282
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 23216 12434 23244 14010
rect 23400 13734 23428 15014
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23124 12406 23244 12434
rect 23308 12434 23336 13330
rect 23492 13190 23520 14894
rect 23584 14890 23612 15914
rect 23726 15260 24022 15280
rect 23782 15258 23806 15260
rect 23862 15258 23886 15260
rect 23942 15258 23966 15260
rect 23804 15206 23806 15258
rect 23868 15206 23880 15258
rect 23942 15206 23944 15258
rect 23782 15204 23806 15206
rect 23862 15204 23886 15206
rect 23942 15204 23966 15206
rect 23726 15184 24022 15204
rect 24216 14952 24268 14958
rect 24214 14920 24216 14929
rect 24268 14920 24270 14929
rect 23572 14884 23624 14890
rect 24214 14855 24270 14864
rect 23572 14826 23624 14832
rect 23584 13784 23612 14826
rect 23726 14172 24022 14192
rect 23782 14170 23806 14172
rect 23862 14170 23886 14172
rect 23942 14170 23966 14172
rect 23804 14118 23806 14170
rect 23868 14118 23880 14170
rect 23942 14118 23944 14170
rect 23782 14116 23806 14118
rect 23862 14116 23886 14118
rect 23942 14116 23966 14118
rect 23726 14096 24022 14116
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 23664 13796 23716 13802
rect 23584 13756 23664 13784
rect 23664 13738 23716 13744
rect 24320 13530 24348 13806
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23726 13084 24022 13104
rect 23782 13082 23806 13084
rect 23862 13082 23886 13084
rect 23942 13082 23966 13084
rect 23804 13030 23806 13082
rect 23868 13030 23880 13082
rect 23942 13030 23944 13082
rect 23782 13028 23806 13030
rect 23862 13028 23886 13030
rect 23942 13028 23966 13030
rect 23726 13008 24022 13028
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23676 12442 23704 12650
rect 23480 12436 23532 12442
rect 23308 12406 23428 12434
rect 23124 11286 23152 12406
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23202 11248 23258 11257
rect 23202 11183 23258 11192
rect 23020 11076 23072 11082
rect 23216 11064 23244 11183
rect 23020 11018 23072 11024
rect 23124 11036 23244 11064
rect 22848 10198 22876 10950
rect 22940 10934 23060 10962
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22940 10198 22968 10406
rect 22836 10192 22888 10198
rect 22836 10134 22888 10140
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 23032 9586 23060 10934
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23124 9518 23152 11036
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22940 8090 22968 9454
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 9042 23060 9318
rect 23216 9178 23244 10474
rect 23308 9586 23336 11494
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 23018 7984 23074 7993
rect 22836 7948 22888 7954
rect 23018 7919 23020 7928
rect 22836 7890 22888 7896
rect 23072 7919 23074 7928
rect 23020 7890 23072 7896
rect 22744 7880 22796 7886
rect 22848 7857 22876 7890
rect 22744 7822 22796 7828
rect 22834 7848 22890 7857
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 6934 22508 7142
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22480 5370 22508 6734
rect 22572 5914 22600 7278
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22664 4146 22692 7278
rect 22756 5914 22784 7822
rect 22834 7783 22890 7792
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22848 7410 22876 7686
rect 23032 7410 23060 7890
rect 22836 7404 22888 7410
rect 23020 7404 23072 7410
rect 22888 7364 22968 7392
rect 22836 7346 22888 7352
rect 22836 7268 22888 7274
rect 22836 7210 22888 7216
rect 22848 6662 22876 7210
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22756 5166 22784 5714
rect 22848 5574 22876 6326
rect 22940 6322 22968 7364
rect 23020 7346 23072 7352
rect 23124 7342 23152 8230
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 23216 6866 23244 8570
rect 23400 7546 23428 12406
rect 23480 12378 23532 12384
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23492 12152 23520 12378
rect 23572 12164 23624 12170
rect 23492 12124 23572 12152
rect 23572 12106 23624 12112
rect 23726 11996 24022 12016
rect 23782 11994 23806 11996
rect 23862 11994 23886 11996
rect 23942 11994 23966 11996
rect 23804 11942 23806 11994
rect 23868 11942 23880 11994
rect 23942 11942 23944 11994
rect 23782 11940 23806 11942
rect 23862 11940 23886 11942
rect 23942 11940 23966 11942
rect 23726 11920 24022 11940
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23492 11354 23520 11630
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23492 10266 23520 11290
rect 23754 11248 23810 11257
rect 24136 11218 24164 13330
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24228 12442 24256 13194
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24412 12306 24440 12582
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24228 11801 24256 12174
rect 24214 11792 24270 11801
rect 24214 11727 24270 11736
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 23754 11183 23756 11192
rect 23808 11183 23810 11192
rect 24124 11212 24176 11218
rect 23756 11154 23808 11160
rect 24124 11154 24176 11160
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 23726 10908 24022 10928
rect 23782 10906 23806 10908
rect 23862 10906 23886 10908
rect 23942 10906 23966 10908
rect 23804 10854 23806 10906
rect 23868 10854 23880 10906
rect 23942 10854 23944 10906
rect 23782 10852 23806 10854
rect 23862 10852 23886 10854
rect 23942 10852 23966 10854
rect 23726 10832 24022 10852
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 24136 10130 24164 10406
rect 24228 10266 24256 11086
rect 24308 11076 24360 11082
rect 24308 11018 24360 11024
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 23584 9382 23612 10066
rect 23726 9820 24022 9840
rect 23782 9818 23806 9820
rect 23862 9818 23886 9820
rect 23942 9818 23966 9820
rect 23804 9766 23806 9818
rect 23868 9766 23880 9818
rect 23942 9766 23944 9818
rect 23782 9764 23806 9766
rect 23862 9764 23886 9766
rect 23942 9764 23966 9766
rect 23726 9744 24022 9764
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 24228 9178 24256 9454
rect 24216 9172 24268 9178
rect 24216 9114 24268 9120
rect 23726 8732 24022 8752
rect 23782 8730 23806 8732
rect 23862 8730 23886 8732
rect 23942 8730 23966 8732
rect 23804 8678 23806 8730
rect 23868 8678 23880 8730
rect 23942 8678 23944 8730
rect 23782 8676 23806 8678
rect 23862 8676 23886 8678
rect 23942 8676 23966 8678
rect 23726 8656 24022 8676
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23492 7546 23520 8366
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 23726 7644 24022 7664
rect 23782 7642 23806 7644
rect 23862 7642 23886 7644
rect 23942 7642 23966 7644
rect 23804 7590 23806 7642
rect 23868 7590 23880 7642
rect 23942 7590 23944 7642
rect 23782 7588 23806 7590
rect 23862 7588 23886 7590
rect 23942 7588 23966 7590
rect 23726 7568 24022 7588
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 23112 6248 23164 6254
rect 23110 6216 23112 6225
rect 23492 6236 23520 7346
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23860 7002 23888 7278
rect 24032 7268 24084 7274
rect 24032 7210 24084 7216
rect 24044 7154 24072 7210
rect 24228 7154 24256 7686
rect 24044 7126 24256 7154
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23584 6730 23704 6746
rect 23584 6724 23716 6730
rect 23584 6718 23664 6724
rect 23584 6458 23612 6718
rect 23664 6666 23716 6672
rect 23726 6556 24022 6576
rect 23782 6554 23806 6556
rect 23862 6554 23886 6556
rect 23942 6554 23966 6556
rect 23804 6502 23806 6554
rect 23868 6502 23880 6554
rect 23942 6502 23944 6554
rect 23782 6500 23806 6502
rect 23862 6500 23886 6502
rect 23942 6500 23966 6502
rect 23726 6480 24022 6500
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23572 6248 23624 6254
rect 23164 6216 23166 6225
rect 23492 6208 23572 6236
rect 23572 6190 23624 6196
rect 23110 6151 23166 6160
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 2122 22692 3878
rect 22756 3670 22784 5102
rect 22848 4622 22876 5306
rect 23032 5166 23060 5646
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 23020 5160 23072 5166
rect 23020 5102 23072 5108
rect 22940 4826 22968 5102
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22744 3664 22796 3670
rect 22744 3606 22796 3612
rect 22848 3058 22876 4558
rect 23032 4457 23060 5102
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23216 4758 23244 4966
rect 23204 4752 23256 4758
rect 23204 4694 23256 4700
rect 23018 4448 23074 4457
rect 23018 4383 23074 4392
rect 23032 3738 23060 4383
rect 23308 4146 23336 6054
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23400 5370 23428 5850
rect 23676 5778 23704 6054
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 23726 5468 24022 5488
rect 23782 5466 23806 5468
rect 23862 5466 23886 5468
rect 23942 5466 23966 5468
rect 23804 5414 23806 5466
rect 23868 5414 23880 5466
rect 23942 5414 23944 5466
rect 23782 5412 23806 5414
rect 23862 5412 23886 5414
rect 23942 5412 23966 5414
rect 23726 5392 24022 5412
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 24136 5098 24164 5510
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 24228 4554 24256 7126
rect 24320 6458 24348 11018
rect 24412 8430 24440 11494
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 24216 4548 24268 4554
rect 24216 4490 24268 4496
rect 23726 4380 24022 4400
rect 23782 4378 23806 4380
rect 23862 4378 23886 4380
rect 23942 4378 23966 4380
rect 23804 4326 23806 4378
rect 23868 4326 23880 4378
rect 23942 4326 23944 4378
rect 23782 4324 23806 4326
rect 23862 4324 23886 4326
rect 23942 4324 23966 4326
rect 23726 4304 24022 4324
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23938 4040 23994 4049
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23216 3398 23244 4014
rect 23400 3942 23428 4014
rect 23938 3975 23940 3984
rect 23992 3975 23994 3984
rect 23940 3946 23992 3952
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23860 3602 23888 3674
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 23216 2582 23244 3334
rect 23400 2650 23428 3538
rect 24320 3534 24348 6190
rect 24400 5840 24452 5846
rect 24400 5782 24452 5788
rect 24412 5370 24440 5782
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24412 3777 24440 4966
rect 24398 3768 24454 3777
rect 24398 3703 24454 3712
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 23726 3292 24022 3312
rect 23782 3290 23806 3292
rect 23862 3290 23886 3292
rect 23942 3290 23966 3292
rect 23804 3238 23806 3290
rect 23868 3238 23880 3290
rect 23942 3238 23944 3290
rect 23782 3236 23806 3238
rect 23862 3236 23886 3238
rect 23942 3236 23966 3238
rect 23726 3216 24022 3236
rect 24136 2990 24164 3334
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 23112 2508 23164 2514
rect 23112 2450 23164 2456
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 22572 2094 22692 2122
rect 22192 1896 22244 1902
rect 22192 1838 22244 1844
rect 21916 1828 21968 1834
rect 21916 1770 21968 1776
rect 22572 800 22600 2094
rect 23032 800 23060 2382
rect 23124 2038 23152 2450
rect 23112 2032 23164 2038
rect 23112 1974 23164 1980
rect 23492 800 23520 2790
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 23726 2204 24022 2224
rect 23782 2202 23806 2204
rect 23862 2202 23886 2204
rect 23942 2202 23966 2204
rect 23804 2150 23806 2202
rect 23868 2150 23880 2202
rect 23942 2150 23944 2202
rect 23782 2148 23806 2150
rect 23862 2148 23886 2150
rect 23942 2148 23966 2150
rect 23726 2128 24022 2148
rect 24136 1970 24164 2246
rect 24124 1964 24176 1970
rect 24124 1906 24176 1912
rect 24412 800 24440 3538
rect 24504 2582 24532 16730
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24596 16114 24624 16390
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24596 13870 24624 14826
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24596 11354 24624 11834
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24596 6458 24624 6802
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24688 6118 24716 27814
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24952 25764 25004 25770
rect 24952 25706 25004 25712
rect 24780 25294 24808 25706
rect 24964 25430 24992 25706
rect 24952 25424 25004 25430
rect 24952 25366 25004 25372
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24780 22250 24808 25230
rect 24780 22222 24900 22250
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 24780 21690 24808 22034
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24872 21570 24900 22222
rect 24780 21542 24900 21570
rect 24780 21418 24808 21542
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24768 20528 24820 20534
rect 24768 20470 24820 20476
rect 24858 20496 24914 20505
rect 24780 18970 24808 20470
rect 24858 20431 24914 20440
rect 24872 20398 24900 20431
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24780 16250 24808 18702
rect 24950 17096 25006 17105
rect 24950 17031 25006 17040
rect 24964 16998 24992 17031
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24872 15162 24900 15914
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24964 14074 24992 15506
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24780 12170 24808 12310
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24780 7750 24808 12106
rect 24872 11898 24900 13330
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24964 11898 24992 12718
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24964 10810 24992 11154
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 25056 9466 25084 28562
rect 25332 28014 25360 30924
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25320 28008 25372 28014
rect 25320 27950 25372 27956
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25240 25430 25268 25638
rect 25228 25424 25280 25430
rect 25228 25366 25280 25372
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25332 22982 25360 23462
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25134 22536 25190 22545
rect 25134 22471 25190 22480
rect 25148 20482 25176 22471
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25424 22234 25452 22374
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25240 21418 25268 22034
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25424 21690 25452 21898
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25608 21570 25636 28970
rect 25792 27606 25820 30924
rect 26146 30696 26202 30705
rect 26146 30631 26202 30640
rect 26054 29336 26110 29345
rect 26054 29271 26110 29280
rect 25964 29096 26016 29102
rect 25964 29038 26016 29044
rect 25976 28014 26004 29038
rect 25964 28008 26016 28014
rect 25964 27950 26016 27956
rect 25780 27600 25832 27606
rect 25780 27542 25832 27548
rect 25780 22500 25832 22506
rect 25780 22442 25832 22448
rect 25792 22234 25820 22442
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25700 21622 25728 22034
rect 25516 21542 25636 21570
rect 25688 21616 25740 21622
rect 25688 21558 25740 21564
rect 25228 21412 25280 21418
rect 25228 21354 25280 21360
rect 25240 21010 25268 21354
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25516 20602 25544 21542
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25608 21010 25636 21422
rect 25700 21350 25728 21558
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25700 21010 25728 21286
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 25792 20856 25820 21286
rect 25700 20828 25820 20856
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25148 20454 25268 20482
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 25148 15745 25176 20266
rect 25240 16402 25268 20454
rect 25700 19417 25728 20828
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25792 19854 25820 20198
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25686 19408 25742 19417
rect 25686 19343 25742 19352
rect 25320 18896 25372 18902
rect 25320 18838 25372 18844
rect 25332 17134 25360 18838
rect 25596 18148 25648 18154
rect 25596 18090 25648 18096
rect 25502 17776 25558 17785
rect 25502 17711 25504 17720
rect 25556 17711 25558 17720
rect 25504 17682 25556 17688
rect 25608 17338 25636 18090
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25240 16374 25360 16402
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25134 15736 25190 15745
rect 25134 15671 25190 15680
rect 25240 14958 25268 16186
rect 25332 16046 25360 16374
rect 25320 16040 25372 16046
rect 25320 15982 25372 15988
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25424 14890 25452 15302
rect 25136 14884 25188 14890
rect 25136 14826 25188 14832
rect 25412 14884 25464 14890
rect 25412 14826 25464 14832
rect 25148 13326 25176 14826
rect 25516 14482 25544 16934
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25608 15745 25636 16594
rect 25594 15736 25650 15745
rect 25594 15671 25650 15680
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25608 14550 25636 15574
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25148 12782 25176 13262
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 24964 9438 25084 9466
rect 25136 9444 25188 9450
rect 24964 9058 24992 9438
rect 25136 9386 25188 9392
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 24872 9030 24992 9058
rect 25056 9042 25084 9318
rect 25044 9036 25096 9042
rect 24872 7954 24900 9030
rect 25044 8978 25096 8984
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24964 8430 24992 8774
rect 25056 8498 25084 8978
rect 25148 8634 25176 9386
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24964 7886 24992 8230
rect 24952 7880 25004 7886
rect 24872 7828 24952 7834
rect 24872 7822 25004 7828
rect 24872 7806 24992 7822
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24872 7342 24900 7806
rect 24964 7757 24992 7806
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 24872 7002 24900 7278
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24766 6216 24822 6225
rect 24766 6151 24822 6160
rect 24780 6118 24808 6151
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24872 5914 24900 6938
rect 25148 6934 25176 8366
rect 25136 6928 25188 6934
rect 25136 6870 25188 6876
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 25240 4570 25268 13466
rect 25424 13462 25452 13942
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25516 12306 25544 12582
rect 25320 12300 25372 12306
rect 25504 12300 25556 12306
rect 25372 12260 25452 12288
rect 25320 12242 25372 12248
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25332 11218 25360 12038
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25424 9058 25452 12260
rect 25504 12242 25556 12248
rect 25516 11694 25544 12242
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25608 11558 25636 14486
rect 25700 14074 25728 19343
rect 25792 19310 25820 19790
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25884 17746 25912 18022
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25792 16658 25820 17614
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25792 13870 25820 14214
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25780 12708 25832 12714
rect 25780 12650 25832 12656
rect 25792 12442 25820 12650
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25608 11286 25636 11494
rect 25596 11280 25648 11286
rect 25596 11222 25648 11228
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 25504 10600 25556 10606
rect 25504 10542 25556 10548
rect 25516 10198 25544 10542
rect 25700 10470 25728 11154
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25792 10606 25820 10950
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25516 9518 25544 10134
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25332 9042 25452 9058
rect 25320 9036 25452 9042
rect 25372 9030 25452 9036
rect 25320 8978 25372 8984
rect 25332 8566 25360 8978
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 6186 25360 7686
rect 25424 6866 25452 8910
rect 25516 8294 25544 9454
rect 25608 9178 25636 10066
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25516 6934 25544 7890
rect 25608 7342 25636 8230
rect 25596 7336 25648 7342
rect 25596 7278 25648 7284
rect 25504 6928 25556 6934
rect 25504 6870 25556 6876
rect 25608 6866 25636 7278
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25320 6180 25372 6186
rect 25320 6122 25372 6128
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 25240 4542 25360 4570
rect 25228 4480 25280 4486
rect 25228 4422 25280 4428
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24780 3194 24808 3470
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 24780 2650 24808 2790
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 24872 800 24900 4014
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24964 2378 24992 3878
rect 25240 3670 25268 4422
rect 25228 3664 25280 3670
rect 25228 3606 25280 3612
rect 25332 2990 25360 4542
rect 25424 3602 25452 4626
rect 25700 3670 25728 10406
rect 25884 8514 25912 16730
rect 25792 8486 25912 8514
rect 25792 8090 25820 8486
rect 25872 8424 25924 8430
rect 25976 8412 26004 27950
rect 26068 27606 26096 29271
rect 26160 29102 26188 30631
rect 26148 29096 26200 29102
rect 26148 29038 26200 29044
rect 26148 28416 26200 28422
rect 26148 28358 26200 28364
rect 26160 27985 26188 28358
rect 26252 28014 26280 30924
rect 27172 29102 27200 30924
rect 27344 29708 27396 29714
rect 27344 29650 27396 29656
rect 27356 29170 27384 29650
rect 27632 29238 27660 30924
rect 28092 29306 28120 30924
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 27620 29232 27672 29238
rect 27620 29174 27672 29180
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27160 29096 27212 29102
rect 27160 29038 27212 29044
rect 26792 29028 26844 29034
rect 26792 28970 26844 28976
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26240 28008 26292 28014
rect 26146 27976 26202 27985
rect 26240 27950 26292 27956
rect 26146 27911 26202 27920
rect 26056 27600 26108 27606
rect 26056 27542 26108 27548
rect 26436 27538 26464 28562
rect 26424 27532 26476 27538
rect 26424 27474 26476 27480
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 26068 24206 26096 25298
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26068 23118 26096 24142
rect 26160 23662 26188 24686
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 23322 26188 23462
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26068 21010 26096 23054
rect 26160 22574 26188 23258
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26252 19334 26280 24550
rect 26344 23497 26372 24618
rect 26436 24410 26464 24618
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26330 23488 26386 23497
rect 26330 23423 26386 23432
rect 26252 19306 26372 19334
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26252 18834 26280 18906
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26252 17814 26280 18566
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26146 17096 26202 17105
rect 26146 17031 26202 17040
rect 26160 16794 26188 17031
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 26056 14884 26108 14890
rect 26056 14826 26108 14832
rect 26068 14346 26096 14826
rect 26146 14376 26202 14385
rect 26056 14340 26108 14346
rect 26146 14311 26202 14320
rect 26056 14282 26108 14288
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 25924 8384 26004 8412
rect 25872 8366 25924 8372
rect 25976 8090 26004 8384
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 26068 7562 26096 14010
rect 26160 14006 26188 14311
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26344 12374 26372 19306
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 26160 11218 26188 11834
rect 26240 11620 26292 11626
rect 26240 11562 26292 11568
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 26252 11150 26280 11562
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 26160 10266 26188 10474
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 26160 9110 26188 10202
rect 26148 9104 26200 9110
rect 26148 9046 26200 9052
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 26252 8022 26280 8502
rect 26240 8016 26292 8022
rect 26240 7958 26292 7964
rect 25884 7534 26096 7562
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 25792 800 25820 3402
rect 25884 2650 25912 7534
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26068 6798 26096 6938
rect 26146 6896 26202 6905
rect 26146 6831 26202 6840
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26160 6254 26188 6831
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 26056 4684 26108 4690
rect 26056 4626 26108 4632
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 25976 1465 26004 4014
rect 25962 1456 26018 1465
rect 25962 1391 26018 1400
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26068 785 26096 4626
rect 26344 4570 26372 11290
rect 26436 9178 26464 23666
rect 26528 22094 26556 27406
rect 26608 25832 26660 25838
rect 26608 25774 26660 25780
rect 26620 25498 26648 25774
rect 26804 25514 26832 28970
rect 29012 28694 29040 30924
rect 29000 28688 29052 28694
rect 26882 28656 26938 28665
rect 29000 28630 29052 28636
rect 26882 28591 26938 28600
rect 26896 27062 26924 28591
rect 27344 27532 27396 27538
rect 27344 27474 27396 27480
rect 26884 27056 26936 27062
rect 26884 26998 26936 27004
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 26882 25936 26938 25945
rect 26882 25871 26884 25880
rect 26936 25871 26938 25880
rect 26884 25842 26936 25848
rect 26608 25492 26660 25498
rect 26804 25486 26924 25514
rect 26608 25434 26660 25440
rect 26608 24744 26660 24750
rect 26608 24686 26660 24692
rect 26620 23662 26648 24686
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 26712 24342 26740 24550
rect 26700 24336 26752 24342
rect 26700 24278 26752 24284
rect 26790 23896 26846 23905
rect 26790 23831 26846 23840
rect 26608 23656 26660 23662
rect 26606 23624 26608 23633
rect 26660 23624 26662 23633
rect 26606 23559 26662 23568
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26712 23254 26740 23462
rect 26700 23248 26752 23254
rect 26700 23190 26752 23196
rect 26804 22574 26832 23831
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26528 22066 26648 22094
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26528 20398 26556 21286
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 26620 19802 26648 22066
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26528 19774 26648 19802
rect 26528 16250 26556 19774
rect 26700 19712 26752 19718
rect 26620 19660 26700 19666
rect 26620 19654 26752 19660
rect 26620 19638 26740 19654
rect 26620 18834 26648 19638
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26620 16726 26648 18770
rect 26712 17134 26740 19246
rect 26804 18970 26832 19858
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26896 18578 26924 25486
rect 26988 25265 27016 26250
rect 27172 25362 27200 26386
rect 27160 25356 27212 25362
rect 27160 25298 27212 25304
rect 26974 25256 27030 25265
rect 26974 25191 27030 25200
rect 26974 23216 27030 23225
rect 26974 23151 27030 23160
rect 26988 22098 27016 23151
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26976 21412 27028 21418
rect 26976 21354 27028 21360
rect 26988 20262 27016 21354
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26988 19938 27016 20198
rect 27080 20058 27108 20946
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 26988 19910 27108 19938
rect 26976 18896 27028 18902
rect 26976 18838 27028 18844
rect 26804 18550 26924 18578
rect 26804 17882 26832 18550
rect 26882 18456 26938 18465
rect 26882 18391 26938 18400
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26896 17270 26924 18391
rect 26988 17542 27016 18838
rect 27080 18426 27108 19910
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 27080 17354 27108 18362
rect 26988 17326 27108 17354
rect 26884 17264 26936 17270
rect 26884 17206 26936 17212
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26608 16720 26660 16726
rect 26608 16662 26660 16668
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26884 15972 26936 15978
rect 26884 15914 26936 15920
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26528 13938 26556 15642
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26712 14958 26740 15302
rect 26896 15065 26924 15914
rect 26882 15056 26938 15065
rect 26882 14991 26938 15000
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26988 13394 27016 17326
rect 27068 15564 27120 15570
rect 27068 15506 27120 15512
rect 27080 14278 27108 15506
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26988 12374 27016 13330
rect 26976 12368 27028 12374
rect 26976 12310 27028 12316
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26516 11688 26568 11694
rect 26896 11665 26924 12038
rect 26516 11630 26568 11636
rect 26882 11656 26938 11665
rect 26528 11354 26556 11630
rect 26882 11591 26938 11600
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26344 4542 26464 4570
rect 26332 4480 26384 4486
rect 26332 4422 26384 4428
rect 26344 4282 26372 4422
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 26146 4040 26202 4049
rect 26146 3975 26202 3984
rect 26160 3942 26188 3975
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 26436 3602 26464 4542
rect 26528 3670 26556 11290
rect 26620 11286 26648 11494
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26790 10296 26846 10305
rect 26790 10231 26846 10240
rect 26698 9616 26754 9625
rect 26698 9551 26754 9560
rect 26712 9518 26740 9551
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26804 9042 26832 10231
rect 26792 9036 26844 9042
rect 26792 8978 26844 8984
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 26712 7585 26740 8366
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26698 7576 26754 7585
rect 26698 7511 26754 7520
rect 26896 6662 26924 8230
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 27172 5642 27200 25298
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27264 15706 27292 22102
rect 27356 21010 27384 27474
rect 27710 26616 27766 26625
rect 27710 26551 27766 26560
rect 27724 26518 27752 26551
rect 27436 26512 27488 26518
rect 27436 26454 27488 26460
rect 27712 26512 27764 26518
rect 27712 26454 27764 26460
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 27344 20800 27396 20806
rect 27344 20742 27396 20748
rect 27356 19310 27384 20742
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 17202 27384 18022
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27252 15700 27304 15706
rect 27252 15642 27304 15648
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27264 11762 27292 15506
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 26804 4185 26832 4626
rect 26790 4176 26846 4185
rect 26790 4111 26846 4120
rect 26516 3664 26568 3670
rect 26516 3606 26568 3612
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26896 3505 26924 5102
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 26882 3496 26938 3505
rect 26516 3460 26568 3466
rect 26882 3431 26938 3440
rect 26516 3402 26568 3408
rect 26240 2916 26292 2922
rect 26240 2858 26292 2864
rect 26252 800 26280 2858
rect 26528 2145 26556 3402
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26514 2136 26570 2145
rect 26514 2071 26570 2080
rect 26804 1442 26832 2790
rect 27080 2582 27108 3538
rect 27356 2990 27384 17138
rect 27448 15570 27476 26454
rect 27528 22160 27580 22166
rect 27528 22102 27580 22108
rect 27540 21185 27568 22102
rect 27618 21992 27674 22001
rect 27618 21927 27674 21936
rect 27632 21894 27660 21927
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27526 21176 27582 21185
rect 27526 21111 27582 21120
rect 27526 19816 27582 19825
rect 27526 19751 27582 19760
rect 27540 18902 27568 19751
rect 27528 18896 27580 18902
rect 27528 18838 27580 18844
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27448 15162 27476 15506
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 27436 14476 27488 14482
rect 27436 14418 27488 14424
rect 27448 5846 27476 14418
rect 27540 10198 27568 17478
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27540 8945 27568 8978
rect 27526 8936 27582 8945
rect 27526 8871 27582 8880
rect 27436 5840 27488 5846
rect 27436 5782 27488 5788
rect 27632 5234 27660 18566
rect 27802 13016 27858 13025
rect 27802 12951 27858 12960
rect 27710 12336 27766 12345
rect 27710 12271 27712 12280
rect 27764 12271 27766 12280
rect 27712 12242 27764 12248
rect 27816 10198 27844 12951
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 27710 8936 27766 8945
rect 27710 8871 27712 8880
rect 27764 8871 27766 8880
rect 27712 8842 27764 8848
rect 27710 6216 27766 6225
rect 27710 6151 27766 6160
rect 27724 5846 27752 6151
rect 27712 5840 27764 5846
rect 27712 5782 27764 5788
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 27526 4856 27582 4865
rect 27526 4791 27582 4800
rect 27540 4758 27568 4791
rect 27528 4752 27580 4758
rect 27528 4694 27580 4700
rect 27620 4004 27672 4010
rect 27620 3946 27672 3952
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 27068 2576 27120 2582
rect 27068 2518 27120 2524
rect 26712 1414 26832 1442
rect 26712 800 26740 1414
rect 27632 800 27660 3946
rect 28540 2508 28592 2514
rect 28540 2450 28592 2456
rect 28080 2372 28132 2378
rect 28080 2314 28132 2320
rect 28092 800 28120 2314
rect 28552 800 28580 2450
rect 26054 776 26110 785
rect 26054 711 26110 720
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28538 0 28594 800
<< via2 >>
rect 1858 29280 1914 29336
rect 2134 28600 2190 28656
rect 1398 27956 1400 27976
rect 1400 27956 1452 27976
rect 1452 27956 1454 27976
rect 1398 27920 1454 27956
rect 1674 25900 1730 25936
rect 1674 25880 1676 25900
rect 1676 25880 1728 25900
rect 1728 25880 1730 25900
rect 1398 25200 1454 25256
rect 1398 17040 1454 17096
rect 1398 15680 1454 15736
rect 1398 15000 1454 15056
rect 1398 12960 1454 13016
rect 1398 9560 1454 9616
rect 1398 8880 1454 8936
rect 1674 23840 1730 23896
rect 1950 26580 2006 26616
rect 1950 26560 1952 26580
rect 1952 26560 2004 26580
rect 2004 26560 2006 26580
rect 1858 23196 1860 23216
rect 1860 23196 1912 23216
rect 1912 23196 1914 23216
rect 1858 23160 1914 23196
rect 2042 22500 2098 22536
rect 2042 22480 2044 22500
rect 2044 22480 2096 22500
rect 2096 22480 2098 22500
rect 1950 21140 2006 21176
rect 1950 21120 1952 21140
rect 1952 21120 2004 21140
rect 2004 21120 2006 21140
rect 1674 20440 1730 20496
rect 1582 18400 1638 18456
rect 1582 17720 1638 17776
rect 1950 19780 2006 19816
rect 1950 19760 1952 19780
rect 1952 19760 2004 19780
rect 2004 19760 2006 19780
rect 2870 30640 2926 30696
rect 5510 29402 5566 29404
rect 5590 29402 5646 29404
rect 5670 29402 5726 29404
rect 5750 29402 5806 29404
rect 5510 29350 5536 29402
rect 5536 29350 5566 29402
rect 5590 29350 5600 29402
rect 5600 29350 5646 29402
rect 5670 29350 5716 29402
rect 5716 29350 5726 29402
rect 5750 29350 5780 29402
rect 5780 29350 5806 29402
rect 5510 29348 5566 29350
rect 5590 29348 5646 29350
rect 5670 29348 5726 29350
rect 5750 29348 5806 29350
rect 1858 14476 1914 14512
rect 1858 14456 1860 14476
rect 1860 14456 1912 14476
rect 1912 14456 1914 14476
rect 2042 14340 2098 14376
rect 2042 14320 2044 14340
rect 2044 14320 2096 14340
rect 2096 14320 2098 14340
rect 2042 12280 2098 12336
rect 1674 11620 1730 11656
rect 1674 11600 1676 11620
rect 1676 11600 1728 11620
rect 1728 11600 1730 11620
rect 1582 7540 1638 7576
rect 1582 7520 1584 7540
rect 1584 7520 1636 7540
rect 1636 7520 1638 7540
rect 1398 6840 1454 6896
rect 1398 6196 1400 6216
rect 1400 6196 1452 6216
rect 1452 6196 1454 6216
rect 1398 6160 1454 6196
rect 1398 4800 1454 4856
rect 1950 10240 2006 10296
rect 4250 21256 4306 21312
rect 4710 19216 4766 19272
rect 2778 4120 2834 4176
rect 1858 1400 1914 1456
rect 3146 3440 3202 3496
rect 4434 7948 4490 7984
rect 4434 7928 4436 7948
rect 4436 7928 4488 7948
rect 4488 7928 4490 7948
rect 2962 2080 3018 2136
rect 5510 28314 5566 28316
rect 5590 28314 5646 28316
rect 5670 28314 5726 28316
rect 5750 28314 5806 28316
rect 5510 28262 5536 28314
rect 5536 28262 5566 28314
rect 5590 28262 5600 28314
rect 5600 28262 5646 28314
rect 5670 28262 5716 28314
rect 5716 28262 5726 28314
rect 5750 28262 5780 28314
rect 5780 28262 5806 28314
rect 5510 28260 5566 28262
rect 5590 28260 5646 28262
rect 5670 28260 5726 28262
rect 5750 28260 5806 28262
rect 5510 27226 5566 27228
rect 5590 27226 5646 27228
rect 5670 27226 5726 27228
rect 5750 27226 5806 27228
rect 5510 27174 5536 27226
rect 5536 27174 5566 27226
rect 5590 27174 5600 27226
rect 5600 27174 5646 27226
rect 5670 27174 5716 27226
rect 5716 27174 5726 27226
rect 5750 27174 5780 27226
rect 5780 27174 5806 27226
rect 5510 27172 5566 27174
rect 5590 27172 5646 27174
rect 5670 27172 5726 27174
rect 5750 27172 5806 27174
rect 5510 26138 5566 26140
rect 5590 26138 5646 26140
rect 5670 26138 5726 26140
rect 5750 26138 5806 26140
rect 5510 26086 5536 26138
rect 5536 26086 5566 26138
rect 5590 26086 5600 26138
rect 5600 26086 5646 26138
rect 5670 26086 5716 26138
rect 5716 26086 5726 26138
rect 5750 26086 5780 26138
rect 5780 26086 5806 26138
rect 5510 26084 5566 26086
rect 5590 26084 5646 26086
rect 5670 26084 5726 26086
rect 5750 26084 5806 26086
rect 5510 25050 5566 25052
rect 5590 25050 5646 25052
rect 5670 25050 5726 25052
rect 5750 25050 5806 25052
rect 5510 24998 5536 25050
rect 5536 24998 5566 25050
rect 5590 24998 5600 25050
rect 5600 24998 5646 25050
rect 5670 24998 5716 25050
rect 5716 24998 5726 25050
rect 5750 24998 5780 25050
rect 5780 24998 5806 25050
rect 5510 24996 5566 24998
rect 5590 24996 5646 24998
rect 5670 24996 5726 24998
rect 5750 24996 5806 24998
rect 5510 23962 5566 23964
rect 5590 23962 5646 23964
rect 5670 23962 5726 23964
rect 5750 23962 5806 23964
rect 5510 23910 5536 23962
rect 5536 23910 5566 23962
rect 5590 23910 5600 23962
rect 5600 23910 5646 23962
rect 5670 23910 5716 23962
rect 5716 23910 5726 23962
rect 5750 23910 5780 23962
rect 5780 23910 5806 23962
rect 5510 23908 5566 23910
rect 5590 23908 5646 23910
rect 5670 23908 5726 23910
rect 5750 23908 5806 23910
rect 5510 22874 5566 22876
rect 5590 22874 5646 22876
rect 5670 22874 5726 22876
rect 5750 22874 5806 22876
rect 5510 22822 5536 22874
rect 5536 22822 5566 22874
rect 5590 22822 5600 22874
rect 5600 22822 5646 22874
rect 5670 22822 5716 22874
rect 5716 22822 5726 22874
rect 5750 22822 5780 22874
rect 5780 22822 5806 22874
rect 5510 22820 5566 22822
rect 5590 22820 5646 22822
rect 5670 22820 5726 22822
rect 5750 22820 5806 22822
rect 5510 21786 5566 21788
rect 5590 21786 5646 21788
rect 5670 21786 5726 21788
rect 5750 21786 5806 21788
rect 5510 21734 5536 21786
rect 5536 21734 5566 21786
rect 5590 21734 5600 21786
rect 5600 21734 5646 21786
rect 5670 21734 5716 21786
rect 5716 21734 5726 21786
rect 5750 21734 5780 21786
rect 5780 21734 5806 21786
rect 5510 21732 5566 21734
rect 5590 21732 5646 21734
rect 5670 21732 5726 21734
rect 5750 21732 5806 21734
rect 5446 21256 5502 21312
rect 5510 20698 5566 20700
rect 5590 20698 5646 20700
rect 5670 20698 5726 20700
rect 5750 20698 5806 20700
rect 5510 20646 5536 20698
rect 5536 20646 5566 20698
rect 5590 20646 5600 20698
rect 5600 20646 5646 20698
rect 5670 20646 5716 20698
rect 5716 20646 5726 20698
rect 5750 20646 5780 20698
rect 5780 20646 5806 20698
rect 5510 20644 5566 20646
rect 5590 20644 5646 20646
rect 5670 20644 5726 20646
rect 5750 20644 5806 20646
rect 5446 19916 5502 19952
rect 5446 19896 5448 19916
rect 5448 19896 5500 19916
rect 5500 19896 5502 19916
rect 5510 19610 5566 19612
rect 5590 19610 5646 19612
rect 5670 19610 5726 19612
rect 5750 19610 5806 19612
rect 5510 19558 5536 19610
rect 5536 19558 5566 19610
rect 5590 19558 5600 19610
rect 5600 19558 5646 19610
rect 5670 19558 5716 19610
rect 5716 19558 5726 19610
rect 5750 19558 5780 19610
rect 5780 19558 5806 19610
rect 5510 19556 5566 19558
rect 5590 19556 5646 19558
rect 5670 19556 5726 19558
rect 5750 19556 5806 19558
rect 5510 18522 5566 18524
rect 5590 18522 5646 18524
rect 5670 18522 5726 18524
rect 5750 18522 5806 18524
rect 5510 18470 5536 18522
rect 5536 18470 5566 18522
rect 5590 18470 5600 18522
rect 5600 18470 5646 18522
rect 5670 18470 5716 18522
rect 5716 18470 5726 18522
rect 5750 18470 5780 18522
rect 5780 18470 5806 18522
rect 5510 18468 5566 18470
rect 5590 18468 5646 18470
rect 5670 18468 5726 18470
rect 5750 18468 5806 18470
rect 7470 28636 7472 28656
rect 7472 28636 7524 28656
rect 7524 28636 7526 28656
rect 7470 28600 7526 28636
rect 5510 17434 5566 17436
rect 5590 17434 5646 17436
rect 5670 17434 5726 17436
rect 5750 17434 5806 17436
rect 5510 17382 5536 17434
rect 5536 17382 5566 17434
rect 5590 17382 5600 17434
rect 5600 17382 5646 17434
rect 5670 17382 5716 17434
rect 5716 17382 5726 17434
rect 5750 17382 5780 17434
rect 5780 17382 5806 17434
rect 5510 17380 5566 17382
rect 5590 17380 5646 17382
rect 5670 17380 5726 17382
rect 5750 17380 5806 17382
rect 4894 12688 4950 12744
rect 6918 21256 6974 21312
rect 5510 16346 5566 16348
rect 5590 16346 5646 16348
rect 5670 16346 5726 16348
rect 5750 16346 5806 16348
rect 5510 16294 5536 16346
rect 5536 16294 5566 16346
rect 5590 16294 5600 16346
rect 5600 16294 5646 16346
rect 5670 16294 5716 16346
rect 5716 16294 5726 16346
rect 5750 16294 5780 16346
rect 5780 16294 5806 16346
rect 5510 16292 5566 16294
rect 5590 16292 5646 16294
rect 5670 16292 5726 16294
rect 5750 16292 5806 16294
rect 5510 15258 5566 15260
rect 5590 15258 5646 15260
rect 5670 15258 5726 15260
rect 5750 15258 5806 15260
rect 5510 15206 5536 15258
rect 5536 15206 5566 15258
rect 5590 15206 5600 15258
rect 5600 15206 5646 15258
rect 5670 15206 5716 15258
rect 5716 15206 5726 15258
rect 5750 15206 5780 15258
rect 5780 15206 5806 15258
rect 5510 15204 5566 15206
rect 5590 15204 5646 15206
rect 5670 15204 5726 15206
rect 5750 15204 5806 15206
rect 5510 14170 5566 14172
rect 5590 14170 5646 14172
rect 5670 14170 5726 14172
rect 5750 14170 5806 14172
rect 5510 14118 5536 14170
rect 5536 14118 5566 14170
rect 5590 14118 5600 14170
rect 5600 14118 5646 14170
rect 5670 14118 5716 14170
rect 5716 14118 5726 14170
rect 5750 14118 5780 14170
rect 5780 14118 5806 14170
rect 5510 14116 5566 14118
rect 5590 14116 5646 14118
rect 5670 14116 5726 14118
rect 5750 14116 5806 14118
rect 5510 13082 5566 13084
rect 5590 13082 5646 13084
rect 5670 13082 5726 13084
rect 5750 13082 5806 13084
rect 5510 13030 5536 13082
rect 5536 13030 5566 13082
rect 5590 13030 5600 13082
rect 5600 13030 5646 13082
rect 5670 13030 5716 13082
rect 5716 13030 5726 13082
rect 5750 13030 5780 13082
rect 5780 13030 5806 13082
rect 5510 13028 5566 13030
rect 5590 13028 5646 13030
rect 5670 13028 5726 13030
rect 5750 13028 5806 13030
rect 5510 11994 5566 11996
rect 5590 11994 5646 11996
rect 5670 11994 5726 11996
rect 5750 11994 5806 11996
rect 5510 11942 5536 11994
rect 5536 11942 5566 11994
rect 5590 11942 5600 11994
rect 5600 11942 5646 11994
rect 5670 11942 5716 11994
rect 5716 11942 5726 11994
rect 5750 11942 5780 11994
rect 5780 11942 5806 11994
rect 5510 11940 5566 11942
rect 5590 11940 5646 11942
rect 5670 11940 5726 11942
rect 5750 11940 5806 11942
rect 5510 10906 5566 10908
rect 5590 10906 5646 10908
rect 5670 10906 5726 10908
rect 5750 10906 5806 10908
rect 5510 10854 5536 10906
rect 5536 10854 5566 10906
rect 5590 10854 5600 10906
rect 5600 10854 5646 10906
rect 5670 10854 5716 10906
rect 5716 10854 5726 10906
rect 5750 10854 5780 10906
rect 5780 10854 5806 10906
rect 5510 10852 5566 10854
rect 5590 10852 5646 10854
rect 5670 10852 5726 10854
rect 5750 10852 5806 10854
rect 5510 9818 5566 9820
rect 5590 9818 5646 9820
rect 5670 9818 5726 9820
rect 5750 9818 5806 9820
rect 5510 9766 5536 9818
rect 5536 9766 5566 9818
rect 5590 9766 5600 9818
rect 5600 9766 5646 9818
rect 5670 9766 5716 9818
rect 5716 9766 5726 9818
rect 5750 9766 5780 9818
rect 5780 9766 5806 9818
rect 5510 9764 5566 9766
rect 5590 9764 5646 9766
rect 5670 9764 5726 9766
rect 5750 9764 5806 9766
rect 5510 8730 5566 8732
rect 5590 8730 5646 8732
rect 5670 8730 5726 8732
rect 5750 8730 5806 8732
rect 5510 8678 5536 8730
rect 5536 8678 5566 8730
rect 5590 8678 5600 8730
rect 5600 8678 5646 8730
rect 5670 8678 5716 8730
rect 5716 8678 5726 8730
rect 5750 8678 5780 8730
rect 5780 8678 5806 8730
rect 5510 8676 5566 8678
rect 5590 8676 5646 8678
rect 5670 8676 5726 8678
rect 5750 8676 5806 8678
rect 5510 7642 5566 7644
rect 5590 7642 5646 7644
rect 5670 7642 5726 7644
rect 5750 7642 5806 7644
rect 5510 7590 5536 7642
rect 5536 7590 5566 7642
rect 5590 7590 5600 7642
rect 5600 7590 5646 7642
rect 5670 7590 5716 7642
rect 5716 7590 5726 7642
rect 5750 7590 5780 7642
rect 5780 7590 5806 7642
rect 5510 7588 5566 7590
rect 5590 7588 5646 7590
rect 5670 7588 5726 7590
rect 5750 7588 5806 7590
rect 6090 7948 6146 7984
rect 6090 7928 6092 7948
rect 6092 7928 6144 7948
rect 6144 7928 6146 7948
rect 5510 6554 5566 6556
rect 5590 6554 5646 6556
rect 5670 6554 5726 6556
rect 5750 6554 5806 6556
rect 5510 6502 5536 6554
rect 5536 6502 5566 6554
rect 5590 6502 5600 6554
rect 5600 6502 5646 6554
rect 5670 6502 5716 6554
rect 5716 6502 5726 6554
rect 5750 6502 5780 6554
rect 5780 6502 5806 6554
rect 5510 6500 5566 6502
rect 5590 6500 5646 6502
rect 5670 6500 5726 6502
rect 5750 6500 5806 6502
rect 6274 6296 6330 6352
rect 5510 5466 5566 5468
rect 5590 5466 5646 5468
rect 5670 5466 5726 5468
rect 5750 5466 5806 5468
rect 5510 5414 5536 5466
rect 5536 5414 5566 5466
rect 5590 5414 5600 5466
rect 5600 5414 5646 5466
rect 5670 5414 5716 5466
rect 5716 5414 5726 5466
rect 5750 5414 5780 5466
rect 5780 5414 5806 5466
rect 5510 5412 5566 5414
rect 5590 5412 5646 5414
rect 5670 5412 5726 5414
rect 5750 5412 5806 5414
rect 5510 4378 5566 4380
rect 5590 4378 5646 4380
rect 5670 4378 5726 4380
rect 5750 4378 5806 4380
rect 5510 4326 5536 4378
rect 5536 4326 5566 4378
rect 5590 4326 5600 4378
rect 5600 4326 5646 4378
rect 5670 4326 5716 4378
rect 5716 4326 5726 4378
rect 5750 4326 5780 4378
rect 5780 4326 5806 4378
rect 5510 4324 5566 4326
rect 5590 4324 5646 4326
rect 5670 4324 5726 4326
rect 5750 4324 5806 4326
rect 5510 3290 5566 3292
rect 5590 3290 5646 3292
rect 5670 3290 5726 3292
rect 5750 3290 5806 3292
rect 5510 3238 5536 3290
rect 5536 3238 5566 3290
rect 5590 3238 5600 3290
rect 5600 3238 5646 3290
rect 5670 3238 5716 3290
rect 5716 3238 5726 3290
rect 5750 3238 5780 3290
rect 5780 3238 5806 3290
rect 5510 3236 5566 3238
rect 5590 3236 5646 3238
rect 5670 3236 5726 3238
rect 5750 3236 5806 3238
rect 7470 19216 7526 19272
rect 7102 12824 7158 12880
rect 7286 12144 7342 12200
rect 8574 28600 8630 28656
rect 10064 28858 10120 28860
rect 10144 28858 10200 28860
rect 10224 28858 10280 28860
rect 10304 28858 10360 28860
rect 10064 28806 10090 28858
rect 10090 28806 10120 28858
rect 10144 28806 10154 28858
rect 10154 28806 10200 28858
rect 10224 28806 10270 28858
rect 10270 28806 10280 28858
rect 10304 28806 10334 28858
rect 10334 28806 10360 28858
rect 10064 28804 10120 28806
rect 10144 28804 10200 28806
rect 10224 28804 10280 28806
rect 10304 28804 10360 28806
rect 9862 28600 9918 28656
rect 9770 27104 9826 27160
rect 10064 27770 10120 27772
rect 10144 27770 10200 27772
rect 10224 27770 10280 27772
rect 10304 27770 10360 27772
rect 10064 27718 10090 27770
rect 10090 27718 10120 27770
rect 10144 27718 10154 27770
rect 10154 27718 10200 27770
rect 10224 27718 10270 27770
rect 10270 27718 10280 27770
rect 10304 27718 10334 27770
rect 10334 27718 10360 27770
rect 10064 27716 10120 27718
rect 10144 27716 10200 27718
rect 10224 27716 10280 27718
rect 10304 27716 10360 27718
rect 9678 26852 9734 26888
rect 9678 26832 9680 26852
rect 9680 26832 9732 26852
rect 9732 26832 9734 26852
rect 8482 19896 8538 19952
rect 7838 14356 7840 14376
rect 7840 14356 7892 14376
rect 7892 14356 7894 14376
rect 7838 14320 7894 14356
rect 7930 12824 7986 12880
rect 7838 12144 7894 12200
rect 8574 14340 8630 14376
rect 8574 14320 8576 14340
rect 8576 14320 8628 14340
rect 8628 14320 8630 14340
rect 10064 26682 10120 26684
rect 10144 26682 10200 26684
rect 10224 26682 10280 26684
rect 10304 26682 10360 26684
rect 10064 26630 10090 26682
rect 10090 26630 10120 26682
rect 10144 26630 10154 26682
rect 10154 26630 10200 26682
rect 10224 26630 10270 26682
rect 10270 26630 10280 26682
rect 10304 26630 10334 26682
rect 10334 26630 10360 26682
rect 10064 26628 10120 26630
rect 10144 26628 10200 26630
rect 10224 26628 10280 26630
rect 10304 26628 10360 26630
rect 10506 27532 10562 27568
rect 10506 27512 10508 27532
rect 10508 27512 10560 27532
rect 10560 27512 10562 27532
rect 10064 25594 10120 25596
rect 10144 25594 10200 25596
rect 10224 25594 10280 25596
rect 10304 25594 10360 25596
rect 10064 25542 10090 25594
rect 10090 25542 10120 25594
rect 10144 25542 10154 25594
rect 10154 25542 10200 25594
rect 10224 25542 10270 25594
rect 10270 25542 10280 25594
rect 10304 25542 10334 25594
rect 10334 25542 10360 25594
rect 10064 25540 10120 25542
rect 10144 25540 10200 25542
rect 10224 25540 10280 25542
rect 10304 25540 10360 25542
rect 10064 24506 10120 24508
rect 10144 24506 10200 24508
rect 10224 24506 10280 24508
rect 10304 24506 10360 24508
rect 10064 24454 10090 24506
rect 10090 24454 10120 24506
rect 10144 24454 10154 24506
rect 10154 24454 10200 24506
rect 10224 24454 10270 24506
rect 10270 24454 10280 24506
rect 10304 24454 10334 24506
rect 10334 24454 10360 24506
rect 10064 24452 10120 24454
rect 10144 24452 10200 24454
rect 10224 24452 10280 24454
rect 10304 24452 10360 24454
rect 9862 24112 9918 24168
rect 9678 21564 9680 21584
rect 9680 21564 9732 21584
rect 9732 21564 9734 21584
rect 9678 21528 9734 21564
rect 10966 25356 11022 25392
rect 10966 25336 10968 25356
rect 10968 25336 11020 25356
rect 11020 25336 11022 25356
rect 10064 23418 10120 23420
rect 10144 23418 10200 23420
rect 10224 23418 10280 23420
rect 10304 23418 10360 23420
rect 10064 23366 10090 23418
rect 10090 23366 10120 23418
rect 10144 23366 10154 23418
rect 10154 23366 10200 23418
rect 10224 23366 10270 23418
rect 10270 23366 10280 23418
rect 10304 23366 10334 23418
rect 10334 23366 10360 23418
rect 10064 23364 10120 23366
rect 10144 23364 10200 23366
rect 10224 23364 10280 23366
rect 10304 23364 10360 23366
rect 10064 22330 10120 22332
rect 10144 22330 10200 22332
rect 10224 22330 10280 22332
rect 10304 22330 10360 22332
rect 10064 22278 10090 22330
rect 10090 22278 10120 22330
rect 10144 22278 10154 22330
rect 10154 22278 10200 22330
rect 10224 22278 10270 22330
rect 10270 22278 10280 22330
rect 10304 22278 10334 22330
rect 10334 22278 10360 22330
rect 10064 22276 10120 22278
rect 10144 22276 10200 22278
rect 10224 22276 10280 22278
rect 10304 22276 10360 22278
rect 10064 21242 10120 21244
rect 10144 21242 10200 21244
rect 10224 21242 10280 21244
rect 10304 21242 10360 21244
rect 10064 21190 10090 21242
rect 10090 21190 10120 21242
rect 10144 21190 10154 21242
rect 10154 21190 10200 21242
rect 10224 21190 10270 21242
rect 10270 21190 10280 21242
rect 10304 21190 10334 21242
rect 10334 21190 10360 21242
rect 10064 21188 10120 21190
rect 10144 21188 10200 21190
rect 10224 21188 10280 21190
rect 10304 21188 10360 21190
rect 10690 23160 10746 23216
rect 10064 20154 10120 20156
rect 10144 20154 10200 20156
rect 10224 20154 10280 20156
rect 10304 20154 10360 20156
rect 10064 20102 10090 20154
rect 10090 20102 10120 20154
rect 10144 20102 10154 20154
rect 10154 20102 10200 20154
rect 10224 20102 10270 20154
rect 10270 20102 10280 20154
rect 10304 20102 10334 20154
rect 10334 20102 10360 20154
rect 10064 20100 10120 20102
rect 10144 20100 10200 20102
rect 10224 20100 10280 20102
rect 10304 20100 10360 20102
rect 10046 19216 10102 19272
rect 10064 19066 10120 19068
rect 10144 19066 10200 19068
rect 10224 19066 10280 19068
rect 10304 19066 10360 19068
rect 10064 19014 10090 19066
rect 10090 19014 10120 19066
rect 10144 19014 10154 19066
rect 10154 19014 10200 19066
rect 10224 19014 10270 19066
rect 10270 19014 10280 19066
rect 10304 19014 10334 19066
rect 10334 19014 10360 19066
rect 10064 19012 10120 19014
rect 10144 19012 10200 19014
rect 10224 19012 10280 19014
rect 10304 19012 10360 19014
rect 10230 18672 10286 18728
rect 10064 17978 10120 17980
rect 10144 17978 10200 17980
rect 10224 17978 10280 17980
rect 10304 17978 10360 17980
rect 10064 17926 10090 17978
rect 10090 17926 10120 17978
rect 10144 17926 10154 17978
rect 10154 17926 10200 17978
rect 10224 17926 10270 17978
rect 10270 17926 10280 17978
rect 10304 17926 10334 17978
rect 10334 17926 10360 17978
rect 10064 17924 10120 17926
rect 10144 17924 10200 17926
rect 10224 17924 10280 17926
rect 10304 17924 10360 17926
rect 9862 17332 9918 17368
rect 9862 17312 9864 17332
rect 9864 17312 9916 17332
rect 9916 17312 9918 17332
rect 9126 14864 9182 14920
rect 9126 14456 9182 14512
rect 5510 2202 5566 2204
rect 5590 2202 5646 2204
rect 5670 2202 5726 2204
rect 5750 2202 5806 2204
rect 5510 2150 5536 2202
rect 5536 2150 5566 2202
rect 5590 2150 5600 2202
rect 5600 2150 5646 2202
rect 5670 2150 5716 2202
rect 5716 2150 5726 2202
rect 5750 2150 5780 2202
rect 5780 2150 5806 2202
rect 5510 2148 5566 2150
rect 5590 2148 5646 2150
rect 5670 2148 5726 2150
rect 5750 2148 5806 2150
rect 8482 10956 8484 10976
rect 8484 10956 8536 10976
rect 8536 10956 8538 10976
rect 8482 10920 8538 10956
rect 8482 6296 8538 6352
rect 8574 5752 8630 5808
rect 9034 11092 9036 11112
rect 9036 11092 9088 11112
rect 9088 11092 9090 11112
rect 9034 11056 9090 11092
rect 9586 14864 9642 14920
rect 10064 16890 10120 16892
rect 10144 16890 10200 16892
rect 10224 16890 10280 16892
rect 10304 16890 10360 16892
rect 10064 16838 10090 16890
rect 10090 16838 10120 16890
rect 10144 16838 10154 16890
rect 10154 16838 10200 16890
rect 10224 16838 10270 16890
rect 10270 16838 10280 16890
rect 10304 16838 10334 16890
rect 10334 16838 10360 16890
rect 10064 16836 10120 16838
rect 10144 16836 10200 16838
rect 10224 16836 10280 16838
rect 10304 16836 10360 16838
rect 10064 15802 10120 15804
rect 10144 15802 10200 15804
rect 10224 15802 10280 15804
rect 10304 15802 10360 15804
rect 10064 15750 10090 15802
rect 10090 15750 10120 15802
rect 10144 15750 10154 15802
rect 10154 15750 10200 15802
rect 10224 15750 10270 15802
rect 10270 15750 10280 15802
rect 10304 15750 10334 15802
rect 10334 15750 10360 15802
rect 10064 15748 10120 15750
rect 10144 15748 10200 15750
rect 10224 15748 10280 15750
rect 10304 15748 10360 15750
rect 10064 14714 10120 14716
rect 10144 14714 10200 14716
rect 10224 14714 10280 14716
rect 10304 14714 10360 14716
rect 10064 14662 10090 14714
rect 10090 14662 10120 14714
rect 10144 14662 10154 14714
rect 10154 14662 10200 14714
rect 10224 14662 10270 14714
rect 10270 14662 10280 14714
rect 10304 14662 10334 14714
rect 10334 14662 10360 14714
rect 10064 14660 10120 14662
rect 10144 14660 10200 14662
rect 10224 14660 10280 14662
rect 10304 14660 10360 14662
rect 9770 13776 9826 13832
rect 10322 14320 10378 14376
rect 9586 12688 9642 12744
rect 10064 13626 10120 13628
rect 10144 13626 10200 13628
rect 10224 13626 10280 13628
rect 10304 13626 10360 13628
rect 10064 13574 10090 13626
rect 10090 13574 10120 13626
rect 10144 13574 10154 13626
rect 10154 13574 10200 13626
rect 10224 13574 10270 13626
rect 10270 13574 10280 13626
rect 10304 13574 10334 13626
rect 10334 13574 10360 13626
rect 10064 13572 10120 13574
rect 10144 13572 10200 13574
rect 10224 13572 10280 13574
rect 10304 13572 10360 13574
rect 12346 24656 12402 24712
rect 11886 19216 11942 19272
rect 12346 18844 12348 18864
rect 12348 18844 12400 18864
rect 12400 18844 12402 18864
rect 12346 18808 12402 18844
rect 11058 16088 11114 16144
rect 10874 15428 10930 15464
rect 10874 15408 10876 15428
rect 10876 15408 10928 15428
rect 10928 15408 10930 15428
rect 10782 14592 10838 14648
rect 10782 13912 10838 13968
rect 10598 13776 10654 13832
rect 10064 12538 10120 12540
rect 10144 12538 10200 12540
rect 10224 12538 10280 12540
rect 10304 12538 10360 12540
rect 10064 12486 10090 12538
rect 10090 12486 10120 12538
rect 10144 12486 10154 12538
rect 10154 12486 10200 12538
rect 10224 12486 10270 12538
rect 10270 12486 10280 12538
rect 10304 12486 10334 12538
rect 10334 12486 10360 12538
rect 10064 12484 10120 12486
rect 10144 12484 10200 12486
rect 10224 12484 10280 12486
rect 10304 12484 10360 12486
rect 10064 11450 10120 11452
rect 10144 11450 10200 11452
rect 10224 11450 10280 11452
rect 10304 11450 10360 11452
rect 10064 11398 10090 11450
rect 10090 11398 10120 11450
rect 10144 11398 10154 11450
rect 10154 11398 10200 11450
rect 10224 11398 10270 11450
rect 10270 11398 10280 11450
rect 10304 11398 10334 11450
rect 10334 11398 10360 11450
rect 10064 11396 10120 11398
rect 10144 11396 10200 11398
rect 10224 11396 10280 11398
rect 10304 11396 10360 11398
rect 10414 10920 10470 10976
rect 10064 10362 10120 10364
rect 10144 10362 10200 10364
rect 10224 10362 10280 10364
rect 10304 10362 10360 10364
rect 10064 10310 10090 10362
rect 10090 10310 10120 10362
rect 10144 10310 10154 10362
rect 10154 10310 10200 10362
rect 10224 10310 10270 10362
rect 10270 10310 10280 10362
rect 10304 10310 10334 10362
rect 10334 10310 10360 10362
rect 10064 10308 10120 10310
rect 10144 10308 10200 10310
rect 10224 10308 10280 10310
rect 10304 10308 10360 10310
rect 9770 8336 9826 8392
rect 10322 9424 10378 9480
rect 10064 9274 10120 9276
rect 10144 9274 10200 9276
rect 10224 9274 10280 9276
rect 10304 9274 10360 9276
rect 10064 9222 10090 9274
rect 10090 9222 10120 9274
rect 10144 9222 10154 9274
rect 10154 9222 10200 9274
rect 10224 9222 10270 9274
rect 10270 9222 10280 9274
rect 10304 9222 10334 9274
rect 10334 9222 10360 9274
rect 10064 9220 10120 9222
rect 10144 9220 10200 9222
rect 10224 9220 10280 9222
rect 10304 9220 10360 9222
rect 10064 8186 10120 8188
rect 10144 8186 10200 8188
rect 10224 8186 10280 8188
rect 10304 8186 10360 8188
rect 10064 8134 10090 8186
rect 10090 8134 10120 8186
rect 10144 8134 10154 8186
rect 10154 8134 10200 8186
rect 10224 8134 10270 8186
rect 10270 8134 10280 8186
rect 10304 8134 10334 8186
rect 10334 8134 10360 8186
rect 10064 8132 10120 8134
rect 10144 8132 10200 8134
rect 10224 8132 10280 8134
rect 10304 8132 10360 8134
rect 10064 7098 10120 7100
rect 10144 7098 10200 7100
rect 10224 7098 10280 7100
rect 10304 7098 10360 7100
rect 10064 7046 10090 7098
rect 10090 7046 10120 7098
rect 10144 7046 10154 7098
rect 10154 7046 10200 7098
rect 10224 7046 10270 7098
rect 10270 7046 10280 7098
rect 10304 7046 10334 7098
rect 10334 7046 10360 7098
rect 10064 7044 10120 7046
rect 10144 7044 10200 7046
rect 10224 7044 10280 7046
rect 10304 7044 10360 7046
rect 9862 5772 9918 5808
rect 9862 5752 9864 5772
rect 9864 5752 9916 5772
rect 9916 5752 9918 5772
rect 10138 6296 10194 6352
rect 10064 6010 10120 6012
rect 10144 6010 10200 6012
rect 10224 6010 10280 6012
rect 10304 6010 10360 6012
rect 10064 5958 10090 6010
rect 10090 5958 10120 6010
rect 10144 5958 10154 6010
rect 10154 5958 10200 6010
rect 10224 5958 10270 6010
rect 10270 5958 10280 6010
rect 10304 5958 10334 6010
rect 10334 5958 10360 6010
rect 10064 5956 10120 5958
rect 10144 5956 10200 5958
rect 10224 5956 10280 5958
rect 10304 5956 10360 5958
rect 9678 3576 9734 3632
rect 10064 4922 10120 4924
rect 10144 4922 10200 4924
rect 10224 4922 10280 4924
rect 10304 4922 10360 4924
rect 10064 4870 10090 4922
rect 10090 4870 10120 4922
rect 10144 4870 10154 4922
rect 10154 4870 10200 4922
rect 10224 4870 10270 4922
rect 10270 4870 10280 4922
rect 10304 4870 10334 4922
rect 10334 4870 10360 4922
rect 10064 4868 10120 4870
rect 10144 4868 10200 4870
rect 10224 4868 10280 4870
rect 10304 4868 10360 4870
rect 10064 3834 10120 3836
rect 10144 3834 10200 3836
rect 10224 3834 10280 3836
rect 10304 3834 10360 3836
rect 10064 3782 10090 3834
rect 10090 3782 10120 3834
rect 10144 3782 10154 3834
rect 10154 3782 10200 3834
rect 10224 3782 10270 3834
rect 10270 3782 10280 3834
rect 10304 3782 10334 3834
rect 10334 3782 10360 3834
rect 10064 3780 10120 3782
rect 10144 3780 10200 3782
rect 10224 3780 10280 3782
rect 10304 3780 10360 3782
rect 10064 2746 10120 2748
rect 10144 2746 10200 2748
rect 10224 2746 10280 2748
rect 10304 2746 10360 2748
rect 10064 2694 10090 2746
rect 10090 2694 10120 2746
rect 10144 2694 10154 2746
rect 10154 2694 10200 2746
rect 10224 2694 10270 2746
rect 10270 2694 10280 2746
rect 10304 2694 10334 2746
rect 10334 2694 10360 2746
rect 10064 2692 10120 2694
rect 10144 2692 10200 2694
rect 10224 2692 10280 2694
rect 10304 2692 10360 2694
rect 9770 2352 9826 2408
rect 10690 11056 10746 11112
rect 12162 13912 12218 13968
rect 14618 29402 14674 29404
rect 14698 29402 14754 29404
rect 14778 29402 14834 29404
rect 14858 29402 14914 29404
rect 14618 29350 14644 29402
rect 14644 29350 14674 29402
rect 14698 29350 14708 29402
rect 14708 29350 14754 29402
rect 14778 29350 14824 29402
rect 14824 29350 14834 29402
rect 14858 29350 14888 29402
rect 14888 29350 14914 29402
rect 14618 29348 14674 29350
rect 14698 29348 14754 29350
rect 14778 29348 14834 29350
rect 14858 29348 14914 29350
rect 14618 28314 14674 28316
rect 14698 28314 14754 28316
rect 14778 28314 14834 28316
rect 14858 28314 14914 28316
rect 14618 28262 14644 28314
rect 14644 28262 14674 28314
rect 14698 28262 14708 28314
rect 14708 28262 14754 28314
rect 14778 28262 14824 28314
rect 14824 28262 14834 28314
rect 14858 28262 14888 28314
rect 14888 28262 14914 28314
rect 14618 28260 14674 28262
rect 14698 28260 14754 28262
rect 14778 28260 14834 28262
rect 14858 28260 14914 28262
rect 13450 25356 13506 25392
rect 13450 25336 13452 25356
rect 13452 25336 13504 25356
rect 13504 25336 13506 25356
rect 14278 24792 14334 24848
rect 13266 21956 13322 21992
rect 13266 21936 13268 21956
rect 13268 21936 13320 21956
rect 13320 21936 13322 21956
rect 13266 21292 13268 21312
rect 13268 21292 13320 21312
rect 13320 21292 13322 21312
rect 13266 21256 13322 21292
rect 13174 18808 13230 18864
rect 12162 10920 12218 10976
rect 12162 9696 12218 9752
rect 13082 15000 13138 15056
rect 10690 4664 10746 4720
rect 11702 4664 11758 4720
rect 12254 6160 12310 6216
rect 12346 3984 12402 4040
rect 12254 3168 12310 3224
rect 12530 4120 12586 4176
rect 12438 2932 12440 2952
rect 12440 2932 12492 2952
rect 12492 2932 12494 2952
rect 12438 2896 12494 2932
rect 12990 3712 13046 3768
rect 12898 3576 12954 3632
rect 15106 27532 15162 27568
rect 15106 27512 15108 27532
rect 15108 27512 15160 27532
rect 15160 27512 15162 27532
rect 14618 27226 14674 27228
rect 14698 27226 14754 27228
rect 14778 27226 14834 27228
rect 14858 27226 14914 27228
rect 14618 27174 14644 27226
rect 14644 27174 14674 27226
rect 14698 27174 14708 27226
rect 14708 27174 14754 27226
rect 14778 27174 14824 27226
rect 14824 27174 14834 27226
rect 14858 27174 14888 27226
rect 14888 27174 14914 27226
rect 14618 27172 14674 27174
rect 14698 27172 14754 27174
rect 14778 27172 14834 27174
rect 14858 27172 14914 27174
rect 14618 26138 14674 26140
rect 14698 26138 14754 26140
rect 14778 26138 14834 26140
rect 14858 26138 14914 26140
rect 14618 26086 14644 26138
rect 14644 26086 14674 26138
rect 14698 26086 14708 26138
rect 14708 26086 14754 26138
rect 14778 26086 14824 26138
rect 14824 26086 14834 26138
rect 14858 26086 14888 26138
rect 14888 26086 14914 26138
rect 14618 26084 14674 26086
rect 14698 26084 14754 26086
rect 14778 26084 14834 26086
rect 14858 26084 14914 26086
rect 14618 25050 14674 25052
rect 14698 25050 14754 25052
rect 14778 25050 14834 25052
rect 14858 25050 14914 25052
rect 14618 24998 14644 25050
rect 14644 24998 14674 25050
rect 14698 24998 14708 25050
rect 14708 24998 14754 25050
rect 14778 24998 14824 25050
rect 14824 24998 14834 25050
rect 14858 24998 14888 25050
rect 14888 24998 14914 25050
rect 14618 24996 14674 24998
rect 14698 24996 14754 24998
rect 14778 24996 14834 24998
rect 14858 24996 14914 24998
rect 14922 24828 14924 24848
rect 14924 24828 14976 24848
rect 14976 24828 14978 24848
rect 14922 24792 14978 24828
rect 14618 23962 14674 23964
rect 14698 23962 14754 23964
rect 14778 23962 14834 23964
rect 14858 23962 14914 23964
rect 14618 23910 14644 23962
rect 14644 23910 14674 23962
rect 14698 23910 14708 23962
rect 14708 23910 14754 23962
rect 14778 23910 14824 23962
rect 14824 23910 14834 23962
rect 14858 23910 14888 23962
rect 14888 23910 14914 23962
rect 14618 23908 14674 23910
rect 14698 23908 14754 23910
rect 14778 23908 14834 23910
rect 14858 23908 14914 23910
rect 14462 23296 14518 23352
rect 14094 21256 14150 21312
rect 14830 23024 14886 23080
rect 14618 22874 14674 22876
rect 14698 22874 14754 22876
rect 14778 22874 14834 22876
rect 14858 22874 14914 22876
rect 14618 22822 14644 22874
rect 14644 22822 14674 22874
rect 14698 22822 14708 22874
rect 14708 22822 14754 22874
rect 14778 22822 14824 22874
rect 14824 22822 14834 22874
rect 14858 22822 14888 22874
rect 14888 22822 14914 22874
rect 14618 22820 14674 22822
rect 14698 22820 14754 22822
rect 14778 22820 14834 22822
rect 14858 22820 14914 22822
rect 14618 21786 14674 21788
rect 14698 21786 14754 21788
rect 14778 21786 14834 21788
rect 14858 21786 14914 21788
rect 14618 21734 14644 21786
rect 14644 21734 14674 21786
rect 14698 21734 14708 21786
rect 14708 21734 14754 21786
rect 14778 21734 14824 21786
rect 14824 21734 14834 21786
rect 14858 21734 14888 21786
rect 14888 21734 14914 21786
rect 14618 21732 14674 21734
rect 14698 21732 14754 21734
rect 14778 21732 14834 21734
rect 14858 21732 14914 21734
rect 14618 20698 14674 20700
rect 14698 20698 14754 20700
rect 14778 20698 14834 20700
rect 14858 20698 14914 20700
rect 14618 20646 14644 20698
rect 14644 20646 14674 20698
rect 14698 20646 14708 20698
rect 14708 20646 14754 20698
rect 14778 20646 14824 20698
rect 14824 20646 14834 20698
rect 14858 20646 14888 20698
rect 14888 20646 14914 20698
rect 14618 20644 14674 20646
rect 14698 20644 14754 20646
rect 14778 20644 14834 20646
rect 14858 20644 14914 20646
rect 15658 24692 15660 24712
rect 15660 24692 15712 24712
rect 15712 24692 15714 24712
rect 15658 24656 15714 24692
rect 14618 19610 14674 19612
rect 14698 19610 14754 19612
rect 14778 19610 14834 19612
rect 14858 19610 14914 19612
rect 14618 19558 14644 19610
rect 14644 19558 14674 19610
rect 14698 19558 14708 19610
rect 14708 19558 14754 19610
rect 14778 19558 14824 19610
rect 14824 19558 14834 19610
rect 14858 19558 14888 19610
rect 14888 19558 14914 19610
rect 14618 19556 14674 19558
rect 14698 19556 14754 19558
rect 14778 19556 14834 19558
rect 14858 19556 14914 19558
rect 14462 18808 14518 18864
rect 14646 18808 14702 18864
rect 14618 18522 14674 18524
rect 14698 18522 14754 18524
rect 14778 18522 14834 18524
rect 14858 18522 14914 18524
rect 14618 18470 14644 18522
rect 14644 18470 14674 18522
rect 14698 18470 14708 18522
rect 14708 18470 14754 18522
rect 14778 18470 14824 18522
rect 14824 18470 14834 18522
rect 14858 18470 14888 18522
rect 14888 18470 14914 18522
rect 14618 18468 14674 18470
rect 14698 18468 14754 18470
rect 14778 18468 14834 18470
rect 14858 18468 14914 18470
rect 15474 19216 15530 19272
rect 15290 18672 15346 18728
rect 14186 17584 14242 17640
rect 14094 16904 14150 16960
rect 14094 14864 14150 14920
rect 14186 14456 14242 14512
rect 14618 17434 14674 17436
rect 14698 17434 14754 17436
rect 14778 17434 14834 17436
rect 14858 17434 14914 17436
rect 14618 17382 14644 17434
rect 14644 17382 14674 17434
rect 14698 17382 14708 17434
rect 14708 17382 14754 17434
rect 14778 17382 14824 17434
rect 14824 17382 14834 17434
rect 14858 17382 14888 17434
rect 14888 17382 14914 17434
rect 14618 17380 14674 17382
rect 14698 17380 14754 17382
rect 14778 17380 14834 17382
rect 14858 17380 14914 17382
rect 14618 16346 14674 16348
rect 14698 16346 14754 16348
rect 14778 16346 14834 16348
rect 14858 16346 14914 16348
rect 14618 16294 14644 16346
rect 14644 16294 14674 16346
rect 14698 16294 14708 16346
rect 14708 16294 14754 16346
rect 14778 16294 14824 16346
rect 14824 16294 14834 16346
rect 14858 16294 14888 16346
rect 14888 16294 14914 16346
rect 14618 16292 14674 16294
rect 14698 16292 14754 16294
rect 14778 16292 14834 16294
rect 14858 16292 14914 16294
rect 14618 15258 14674 15260
rect 14698 15258 14754 15260
rect 14778 15258 14834 15260
rect 14858 15258 14914 15260
rect 14618 15206 14644 15258
rect 14644 15206 14674 15258
rect 14698 15206 14708 15258
rect 14708 15206 14754 15258
rect 14778 15206 14824 15258
rect 14824 15206 14834 15258
rect 14858 15206 14888 15258
rect 14888 15206 14914 15258
rect 14618 15204 14674 15206
rect 14698 15204 14754 15206
rect 14778 15204 14834 15206
rect 14858 15204 14914 15206
rect 14830 14884 14886 14920
rect 14830 14864 14832 14884
rect 14832 14864 14884 14884
rect 14884 14864 14886 14884
rect 14922 14728 14978 14784
rect 14738 14320 14794 14376
rect 14618 14170 14674 14172
rect 14698 14170 14754 14172
rect 14778 14170 14834 14172
rect 14858 14170 14914 14172
rect 14618 14118 14644 14170
rect 14644 14118 14674 14170
rect 14698 14118 14708 14170
rect 14708 14118 14754 14170
rect 14778 14118 14824 14170
rect 14824 14118 14834 14170
rect 14858 14118 14888 14170
rect 14888 14118 14914 14170
rect 14618 14116 14674 14118
rect 14698 14116 14754 14118
rect 14778 14116 14834 14118
rect 14858 14116 14914 14118
rect 14618 13082 14674 13084
rect 14698 13082 14754 13084
rect 14778 13082 14834 13084
rect 14858 13082 14914 13084
rect 14618 13030 14644 13082
rect 14644 13030 14674 13082
rect 14698 13030 14708 13082
rect 14708 13030 14754 13082
rect 14778 13030 14824 13082
rect 14824 13030 14834 13082
rect 14858 13030 14888 13082
rect 14888 13030 14914 13082
rect 14618 13028 14674 13030
rect 14698 13028 14754 13030
rect 14778 13028 14834 13030
rect 14858 13028 14914 13030
rect 13542 8356 13598 8392
rect 13542 8336 13544 8356
rect 13544 8336 13596 8356
rect 13596 8336 13598 8356
rect 13266 4684 13322 4720
rect 13266 4664 13268 4684
rect 13268 4664 13320 4684
rect 13320 4664 13322 4684
rect 13174 3984 13230 4040
rect 12898 3168 12954 3224
rect 13910 9696 13966 9752
rect 15198 16244 15254 16280
rect 15198 16224 15200 16244
rect 15200 16224 15252 16244
rect 15252 16224 15254 16244
rect 15198 14728 15254 14784
rect 14618 11994 14674 11996
rect 14698 11994 14754 11996
rect 14778 11994 14834 11996
rect 14858 11994 14914 11996
rect 14618 11942 14644 11994
rect 14644 11942 14674 11994
rect 14698 11942 14708 11994
rect 14708 11942 14754 11994
rect 14778 11942 14824 11994
rect 14824 11942 14834 11994
rect 14858 11942 14888 11994
rect 14888 11942 14914 11994
rect 14618 11940 14674 11942
rect 14698 11940 14754 11942
rect 14778 11940 14834 11942
rect 14858 11940 14914 11942
rect 15566 14864 15622 14920
rect 15934 24792 15990 24848
rect 16026 16904 16082 16960
rect 15934 16124 15936 16144
rect 15936 16124 15988 16144
rect 15988 16124 15990 16144
rect 15934 16088 15990 16124
rect 14618 10906 14674 10908
rect 14698 10906 14754 10908
rect 14778 10906 14834 10908
rect 14858 10906 14914 10908
rect 14618 10854 14644 10906
rect 14644 10854 14674 10906
rect 14698 10854 14708 10906
rect 14708 10854 14754 10906
rect 14778 10854 14824 10906
rect 14824 10854 14834 10906
rect 14858 10854 14888 10906
rect 14888 10854 14914 10906
rect 14618 10852 14674 10854
rect 14698 10852 14754 10854
rect 14778 10852 14834 10854
rect 14858 10852 14914 10854
rect 14618 9818 14674 9820
rect 14698 9818 14754 9820
rect 14778 9818 14834 9820
rect 14858 9818 14914 9820
rect 14618 9766 14644 9818
rect 14644 9766 14674 9818
rect 14698 9766 14708 9818
rect 14708 9766 14754 9818
rect 14778 9766 14824 9818
rect 14824 9766 14834 9818
rect 14858 9766 14888 9818
rect 14888 9766 14914 9818
rect 14618 9764 14674 9766
rect 14698 9764 14754 9766
rect 14778 9764 14834 9766
rect 14858 9764 14914 9766
rect 14618 8730 14674 8732
rect 14698 8730 14754 8732
rect 14778 8730 14834 8732
rect 14858 8730 14914 8732
rect 14618 8678 14644 8730
rect 14644 8678 14674 8730
rect 14698 8678 14708 8730
rect 14708 8678 14754 8730
rect 14778 8678 14824 8730
rect 14824 8678 14834 8730
rect 14858 8678 14888 8730
rect 14888 8678 14914 8730
rect 14618 8676 14674 8678
rect 14698 8676 14754 8678
rect 14778 8676 14834 8678
rect 14858 8676 14914 8678
rect 14186 8472 14242 8528
rect 16302 15408 16358 15464
rect 15750 12824 15806 12880
rect 15934 12552 15990 12608
rect 15842 12416 15898 12472
rect 16210 13776 16266 13832
rect 14618 7642 14674 7644
rect 14698 7642 14754 7644
rect 14778 7642 14834 7644
rect 14858 7642 14914 7644
rect 14618 7590 14644 7642
rect 14644 7590 14674 7642
rect 14698 7590 14708 7642
rect 14708 7590 14754 7642
rect 14778 7590 14824 7642
rect 14824 7590 14834 7642
rect 14858 7590 14888 7642
rect 14888 7590 14914 7642
rect 14618 7588 14674 7590
rect 14698 7588 14754 7590
rect 14778 7588 14834 7590
rect 14858 7588 14914 7590
rect 14618 6554 14674 6556
rect 14698 6554 14754 6556
rect 14778 6554 14834 6556
rect 14858 6554 14914 6556
rect 14618 6502 14644 6554
rect 14644 6502 14674 6554
rect 14698 6502 14708 6554
rect 14708 6502 14754 6554
rect 14778 6502 14824 6554
rect 14824 6502 14834 6554
rect 14858 6502 14888 6554
rect 14888 6502 14914 6554
rect 14618 6500 14674 6502
rect 14698 6500 14754 6502
rect 14778 6500 14834 6502
rect 14858 6500 14914 6502
rect 14002 6196 14004 6216
rect 14004 6196 14056 6216
rect 14056 6196 14058 6216
rect 14002 6160 14058 6196
rect 14618 5466 14674 5468
rect 14698 5466 14754 5468
rect 14778 5466 14834 5468
rect 14858 5466 14914 5468
rect 14618 5414 14644 5466
rect 14644 5414 14674 5466
rect 14698 5414 14708 5466
rect 14708 5414 14754 5466
rect 14778 5414 14824 5466
rect 14824 5414 14834 5466
rect 14858 5414 14888 5466
rect 14888 5414 14914 5466
rect 14618 5412 14674 5414
rect 14698 5412 14754 5414
rect 14778 5412 14834 5414
rect 14858 5412 14914 5414
rect 14618 4378 14674 4380
rect 14698 4378 14754 4380
rect 14778 4378 14834 4380
rect 14858 4378 14914 4380
rect 14618 4326 14644 4378
rect 14644 4326 14674 4378
rect 14698 4326 14708 4378
rect 14708 4326 14754 4378
rect 14778 4326 14824 4378
rect 14824 4326 14834 4378
rect 14858 4326 14888 4378
rect 14888 4326 14914 4378
rect 14618 4324 14674 4326
rect 14698 4324 14754 4326
rect 14778 4324 14834 4326
rect 14858 4324 14914 4326
rect 14618 3290 14674 3292
rect 14698 3290 14754 3292
rect 14778 3290 14834 3292
rect 14858 3290 14914 3292
rect 14618 3238 14644 3290
rect 14644 3238 14674 3290
rect 14698 3238 14708 3290
rect 14708 3238 14754 3290
rect 14778 3238 14824 3290
rect 14824 3238 14834 3290
rect 14858 3238 14888 3290
rect 14888 3238 14914 3290
rect 14618 3236 14674 3238
rect 14698 3236 14754 3238
rect 14778 3236 14834 3238
rect 14858 3236 14914 3238
rect 14618 2202 14674 2204
rect 14698 2202 14754 2204
rect 14778 2202 14834 2204
rect 14858 2202 14914 2204
rect 14618 2150 14644 2202
rect 14644 2150 14674 2202
rect 14698 2150 14708 2202
rect 14708 2150 14754 2202
rect 14778 2150 14824 2202
rect 14824 2150 14834 2202
rect 14858 2150 14888 2202
rect 14888 2150 14914 2202
rect 14618 2148 14674 2150
rect 14698 2148 14754 2150
rect 14778 2148 14834 2150
rect 14858 2148 14914 2150
rect 15474 3460 15530 3496
rect 15474 3440 15476 3460
rect 15476 3440 15528 3460
rect 15528 3440 15530 3460
rect 16670 17604 16726 17640
rect 16670 17584 16672 17604
rect 16672 17584 16724 17604
rect 16724 17584 16726 17604
rect 19172 28858 19228 28860
rect 19252 28858 19308 28860
rect 19332 28858 19388 28860
rect 19412 28858 19468 28860
rect 19172 28806 19198 28858
rect 19198 28806 19228 28858
rect 19252 28806 19262 28858
rect 19262 28806 19308 28858
rect 19332 28806 19378 28858
rect 19378 28806 19388 28858
rect 19412 28806 19442 28858
rect 19442 28806 19468 28858
rect 19172 28804 19228 28806
rect 19252 28804 19308 28806
rect 19332 28804 19388 28806
rect 19412 28804 19468 28806
rect 19172 27770 19228 27772
rect 19252 27770 19308 27772
rect 19332 27770 19388 27772
rect 19412 27770 19468 27772
rect 19172 27718 19198 27770
rect 19198 27718 19228 27770
rect 19252 27718 19262 27770
rect 19262 27718 19308 27770
rect 19332 27718 19378 27770
rect 19378 27718 19388 27770
rect 19412 27718 19442 27770
rect 19442 27718 19468 27770
rect 19172 27716 19228 27718
rect 19252 27716 19308 27718
rect 19332 27716 19388 27718
rect 19412 27716 19468 27718
rect 17130 18672 17186 18728
rect 17222 14476 17278 14512
rect 17222 14456 17224 14476
rect 17224 14456 17276 14476
rect 17276 14456 17278 14476
rect 16854 11872 16910 11928
rect 16118 3984 16174 4040
rect 17590 18672 17646 18728
rect 17590 14592 17646 14648
rect 17314 11872 17370 11928
rect 16302 3032 16358 3088
rect 16670 2896 16726 2952
rect 17222 4392 17278 4448
rect 18050 16940 18052 16960
rect 18052 16940 18104 16960
rect 18104 16940 18106 16960
rect 18050 16904 18106 16940
rect 17958 14592 18014 14648
rect 17958 13912 18014 13968
rect 18234 22072 18290 22128
rect 18234 21528 18290 21584
rect 18234 21428 18236 21448
rect 18236 21428 18288 21448
rect 18288 21428 18290 21448
rect 18234 21392 18290 21428
rect 19172 26682 19228 26684
rect 19252 26682 19308 26684
rect 19332 26682 19388 26684
rect 19412 26682 19468 26684
rect 19172 26630 19198 26682
rect 19198 26630 19228 26682
rect 19252 26630 19262 26682
rect 19262 26630 19308 26682
rect 19332 26630 19378 26682
rect 19378 26630 19388 26682
rect 19412 26630 19442 26682
rect 19442 26630 19468 26682
rect 19172 26628 19228 26630
rect 19252 26628 19308 26630
rect 19332 26628 19388 26630
rect 19412 26628 19468 26630
rect 19172 25594 19228 25596
rect 19252 25594 19308 25596
rect 19332 25594 19388 25596
rect 19412 25594 19468 25596
rect 19172 25542 19198 25594
rect 19198 25542 19228 25594
rect 19252 25542 19262 25594
rect 19262 25542 19308 25594
rect 19332 25542 19378 25594
rect 19378 25542 19388 25594
rect 19412 25542 19442 25594
rect 19442 25542 19468 25594
rect 19172 25540 19228 25542
rect 19252 25540 19308 25542
rect 19332 25540 19388 25542
rect 19412 25540 19468 25542
rect 18786 23296 18842 23352
rect 18694 23160 18750 23216
rect 18234 16224 18290 16280
rect 18234 13912 18290 13968
rect 18234 12824 18290 12880
rect 18510 14728 18566 14784
rect 18510 14476 18566 14512
rect 18510 14456 18512 14476
rect 18512 14456 18564 14476
rect 18564 14456 18566 14476
rect 18326 12552 18382 12608
rect 17682 6296 17738 6352
rect 19172 24506 19228 24508
rect 19252 24506 19308 24508
rect 19332 24506 19388 24508
rect 19412 24506 19468 24508
rect 19172 24454 19198 24506
rect 19198 24454 19228 24506
rect 19252 24454 19262 24506
rect 19262 24454 19308 24506
rect 19332 24454 19378 24506
rect 19378 24454 19388 24506
rect 19412 24454 19442 24506
rect 19442 24454 19468 24506
rect 19172 24452 19228 24454
rect 19252 24452 19308 24454
rect 19332 24452 19388 24454
rect 19412 24452 19468 24454
rect 19172 23418 19228 23420
rect 19252 23418 19308 23420
rect 19332 23418 19388 23420
rect 19412 23418 19468 23420
rect 19172 23366 19198 23418
rect 19198 23366 19228 23418
rect 19252 23366 19262 23418
rect 19262 23366 19308 23418
rect 19332 23366 19378 23418
rect 19378 23366 19388 23418
rect 19412 23366 19442 23418
rect 19442 23366 19468 23418
rect 19172 23364 19228 23366
rect 19252 23364 19308 23366
rect 19332 23364 19388 23366
rect 19412 23364 19468 23366
rect 19154 23024 19210 23080
rect 19172 22330 19228 22332
rect 19252 22330 19308 22332
rect 19332 22330 19388 22332
rect 19412 22330 19468 22332
rect 19172 22278 19198 22330
rect 19198 22278 19228 22330
rect 19252 22278 19262 22330
rect 19262 22278 19308 22330
rect 19332 22278 19378 22330
rect 19378 22278 19388 22330
rect 19412 22278 19442 22330
rect 19442 22278 19468 22330
rect 19172 22276 19228 22278
rect 19252 22276 19308 22278
rect 19332 22276 19388 22278
rect 19412 22276 19468 22278
rect 19246 21392 19302 21448
rect 19172 21242 19228 21244
rect 19252 21242 19308 21244
rect 19332 21242 19388 21244
rect 19412 21242 19468 21244
rect 19172 21190 19198 21242
rect 19198 21190 19228 21242
rect 19252 21190 19262 21242
rect 19262 21190 19308 21242
rect 19332 21190 19378 21242
rect 19378 21190 19388 21242
rect 19412 21190 19442 21242
rect 19442 21190 19468 21242
rect 19172 21188 19228 21190
rect 19252 21188 19308 21190
rect 19332 21188 19388 21190
rect 19412 21188 19468 21190
rect 19172 20154 19228 20156
rect 19252 20154 19308 20156
rect 19332 20154 19388 20156
rect 19412 20154 19468 20156
rect 19172 20102 19198 20154
rect 19198 20102 19228 20154
rect 19252 20102 19262 20154
rect 19262 20102 19308 20154
rect 19332 20102 19378 20154
rect 19378 20102 19388 20154
rect 19412 20102 19442 20154
rect 19442 20102 19468 20154
rect 19172 20100 19228 20102
rect 19252 20100 19308 20102
rect 19332 20100 19388 20102
rect 19412 20100 19468 20102
rect 19172 19066 19228 19068
rect 19252 19066 19308 19068
rect 19332 19066 19388 19068
rect 19412 19066 19468 19068
rect 19172 19014 19198 19066
rect 19198 19014 19228 19066
rect 19252 19014 19262 19066
rect 19262 19014 19308 19066
rect 19332 19014 19378 19066
rect 19378 19014 19388 19066
rect 19412 19014 19442 19066
rect 19442 19014 19468 19066
rect 19172 19012 19228 19014
rect 19252 19012 19308 19014
rect 19332 19012 19388 19014
rect 19412 19012 19468 19014
rect 18510 3440 18566 3496
rect 18970 15000 19026 15056
rect 19172 17978 19228 17980
rect 19252 17978 19308 17980
rect 19332 17978 19388 17980
rect 19412 17978 19468 17980
rect 19172 17926 19198 17978
rect 19198 17926 19228 17978
rect 19252 17926 19262 17978
rect 19262 17926 19308 17978
rect 19332 17926 19378 17978
rect 19378 17926 19388 17978
rect 19412 17926 19442 17978
rect 19442 17926 19468 17978
rect 19172 17924 19228 17926
rect 19252 17924 19308 17926
rect 19332 17924 19388 17926
rect 19412 17924 19468 17926
rect 19614 17196 19670 17232
rect 19614 17176 19616 17196
rect 19616 17176 19668 17196
rect 19668 17176 19670 17196
rect 19172 16890 19228 16892
rect 19252 16890 19308 16892
rect 19332 16890 19388 16892
rect 19412 16890 19468 16892
rect 19172 16838 19198 16890
rect 19198 16838 19228 16890
rect 19252 16838 19262 16890
rect 19262 16838 19308 16890
rect 19332 16838 19378 16890
rect 19378 16838 19388 16890
rect 19412 16838 19442 16890
rect 19442 16838 19468 16890
rect 19172 16836 19228 16838
rect 19252 16836 19308 16838
rect 19332 16836 19388 16838
rect 19412 16836 19468 16838
rect 19982 19352 20038 19408
rect 19982 18164 19984 18184
rect 19984 18164 20036 18184
rect 20036 18164 20038 18184
rect 19982 18128 20038 18164
rect 19172 15802 19228 15804
rect 19252 15802 19308 15804
rect 19332 15802 19388 15804
rect 19412 15802 19468 15804
rect 19172 15750 19198 15802
rect 19198 15750 19228 15802
rect 19252 15750 19262 15802
rect 19262 15750 19308 15802
rect 19332 15750 19378 15802
rect 19378 15750 19388 15802
rect 19412 15750 19442 15802
rect 19442 15750 19468 15802
rect 19172 15748 19228 15750
rect 19252 15748 19308 15750
rect 19332 15748 19388 15750
rect 19412 15748 19468 15750
rect 19172 14714 19228 14716
rect 19252 14714 19308 14716
rect 19332 14714 19388 14716
rect 19412 14714 19468 14716
rect 19172 14662 19198 14714
rect 19198 14662 19228 14714
rect 19252 14662 19262 14714
rect 19262 14662 19308 14714
rect 19332 14662 19378 14714
rect 19378 14662 19388 14714
rect 19412 14662 19442 14714
rect 19442 14662 19468 14714
rect 19172 14660 19228 14662
rect 19252 14660 19308 14662
rect 19332 14660 19388 14662
rect 19412 14660 19468 14662
rect 19172 13626 19228 13628
rect 19252 13626 19308 13628
rect 19332 13626 19388 13628
rect 19412 13626 19468 13628
rect 19172 13574 19198 13626
rect 19198 13574 19228 13626
rect 19252 13574 19262 13626
rect 19262 13574 19308 13626
rect 19332 13574 19378 13626
rect 19378 13574 19388 13626
rect 19412 13574 19442 13626
rect 19442 13574 19468 13626
rect 19172 13572 19228 13574
rect 19252 13572 19308 13574
rect 19332 13572 19388 13574
rect 19412 13572 19468 13574
rect 18970 12416 19026 12472
rect 19172 12538 19228 12540
rect 19252 12538 19308 12540
rect 19332 12538 19388 12540
rect 19412 12538 19468 12540
rect 19172 12486 19198 12538
rect 19198 12486 19228 12538
rect 19252 12486 19262 12538
rect 19262 12486 19308 12538
rect 19332 12486 19378 12538
rect 19378 12486 19388 12538
rect 19412 12486 19442 12538
rect 19442 12486 19468 12538
rect 19172 12484 19228 12486
rect 19252 12484 19308 12486
rect 19332 12484 19388 12486
rect 19412 12484 19468 12486
rect 19172 11450 19228 11452
rect 19252 11450 19308 11452
rect 19332 11450 19388 11452
rect 19412 11450 19468 11452
rect 19172 11398 19198 11450
rect 19198 11398 19228 11450
rect 19252 11398 19262 11450
rect 19262 11398 19308 11450
rect 19332 11398 19378 11450
rect 19378 11398 19388 11450
rect 19412 11398 19442 11450
rect 19442 11398 19468 11450
rect 19172 11396 19228 11398
rect 19252 11396 19308 11398
rect 19332 11396 19388 11398
rect 19412 11396 19468 11398
rect 19172 10362 19228 10364
rect 19252 10362 19308 10364
rect 19332 10362 19388 10364
rect 19412 10362 19468 10364
rect 19172 10310 19198 10362
rect 19198 10310 19228 10362
rect 19252 10310 19262 10362
rect 19262 10310 19308 10362
rect 19332 10310 19378 10362
rect 19378 10310 19388 10362
rect 19412 10310 19442 10362
rect 19442 10310 19468 10362
rect 19172 10308 19228 10310
rect 19252 10308 19308 10310
rect 19332 10308 19388 10310
rect 19412 10308 19468 10310
rect 19890 15272 19946 15328
rect 19706 14864 19762 14920
rect 19172 9274 19228 9276
rect 19252 9274 19308 9276
rect 19332 9274 19388 9276
rect 19412 9274 19468 9276
rect 19172 9222 19198 9274
rect 19198 9222 19228 9274
rect 19252 9222 19262 9274
rect 19262 9222 19308 9274
rect 19332 9222 19378 9274
rect 19378 9222 19388 9274
rect 19412 9222 19442 9274
rect 19442 9222 19468 9274
rect 19172 9220 19228 9222
rect 19252 9220 19308 9222
rect 19332 9220 19388 9222
rect 19412 9220 19468 9222
rect 19890 8916 19892 8936
rect 19892 8916 19944 8936
rect 19944 8916 19946 8936
rect 19890 8880 19946 8916
rect 18970 8472 19026 8528
rect 19172 8186 19228 8188
rect 19252 8186 19308 8188
rect 19332 8186 19388 8188
rect 19412 8186 19468 8188
rect 19172 8134 19198 8186
rect 19198 8134 19228 8186
rect 19252 8134 19262 8186
rect 19262 8134 19308 8186
rect 19332 8134 19378 8186
rect 19378 8134 19388 8186
rect 19412 8134 19442 8186
rect 19442 8134 19468 8186
rect 19172 8132 19228 8134
rect 19252 8132 19308 8134
rect 19332 8132 19388 8134
rect 19412 8132 19468 8134
rect 20718 17040 20774 17096
rect 20902 22072 20958 22128
rect 20994 18128 21050 18184
rect 23726 29402 23782 29404
rect 23806 29402 23862 29404
rect 23886 29402 23942 29404
rect 23966 29402 24022 29404
rect 23726 29350 23752 29402
rect 23752 29350 23782 29402
rect 23806 29350 23816 29402
rect 23816 29350 23862 29402
rect 23886 29350 23932 29402
rect 23932 29350 23942 29402
rect 23966 29350 23996 29402
rect 23996 29350 24022 29402
rect 23726 29348 23782 29350
rect 23806 29348 23862 29350
rect 23886 29348 23942 29350
rect 23966 29348 24022 29350
rect 21270 23568 21326 23624
rect 21546 17176 21602 17232
rect 20810 15680 20866 15736
rect 20810 11736 20866 11792
rect 21362 14884 21418 14920
rect 21362 14864 21364 14884
rect 21364 14864 21416 14884
rect 21416 14864 21418 14884
rect 20902 9560 20958 9616
rect 21178 11736 21234 11792
rect 21270 11192 21326 11248
rect 20902 7948 20958 7984
rect 20902 7928 20904 7948
rect 20904 7928 20956 7948
rect 20956 7928 20958 7948
rect 20258 7792 20314 7848
rect 19172 7098 19228 7100
rect 19252 7098 19308 7100
rect 19332 7098 19388 7100
rect 19412 7098 19468 7100
rect 19172 7046 19198 7098
rect 19198 7046 19228 7098
rect 19252 7046 19262 7098
rect 19262 7046 19308 7098
rect 19332 7046 19378 7098
rect 19378 7046 19388 7098
rect 19412 7046 19442 7098
rect 19442 7046 19468 7098
rect 19172 7044 19228 7046
rect 19252 7044 19308 7046
rect 19332 7044 19388 7046
rect 19412 7044 19468 7046
rect 19172 6010 19228 6012
rect 19252 6010 19308 6012
rect 19332 6010 19388 6012
rect 19412 6010 19468 6012
rect 19172 5958 19198 6010
rect 19198 5958 19228 6010
rect 19252 5958 19262 6010
rect 19262 5958 19308 6010
rect 19332 5958 19378 6010
rect 19378 5958 19388 6010
rect 19412 5958 19442 6010
rect 19442 5958 19468 6010
rect 19172 5956 19228 5958
rect 19252 5956 19308 5958
rect 19332 5956 19388 5958
rect 19412 5956 19468 5958
rect 19172 4922 19228 4924
rect 19252 4922 19308 4924
rect 19332 4922 19388 4924
rect 19412 4922 19468 4924
rect 19172 4870 19198 4922
rect 19198 4870 19228 4922
rect 19252 4870 19262 4922
rect 19262 4870 19308 4922
rect 19332 4870 19378 4922
rect 19378 4870 19388 4922
rect 19412 4870 19442 4922
rect 19442 4870 19468 4922
rect 19172 4868 19228 4870
rect 19252 4868 19308 4870
rect 19332 4868 19388 4870
rect 19412 4868 19468 4870
rect 19172 3834 19228 3836
rect 19252 3834 19308 3836
rect 19332 3834 19388 3836
rect 19412 3834 19468 3836
rect 19172 3782 19198 3834
rect 19198 3782 19228 3834
rect 19252 3782 19262 3834
rect 19262 3782 19308 3834
rect 19332 3782 19378 3834
rect 19378 3782 19388 3834
rect 19412 3782 19442 3834
rect 19442 3782 19468 3834
rect 19172 3780 19228 3782
rect 19252 3780 19308 3782
rect 19332 3780 19388 3782
rect 19412 3780 19468 3782
rect 19154 3576 19210 3632
rect 19338 2896 19394 2952
rect 19172 2746 19228 2748
rect 19252 2746 19308 2748
rect 19332 2746 19388 2748
rect 19412 2746 19468 2748
rect 19172 2694 19198 2746
rect 19198 2694 19228 2746
rect 19252 2694 19262 2746
rect 19262 2694 19308 2746
rect 19332 2694 19378 2746
rect 19378 2694 19388 2746
rect 19412 2694 19442 2746
rect 19442 2694 19468 2746
rect 19172 2692 19228 2694
rect 19252 2692 19308 2694
rect 19332 2692 19388 2694
rect 19412 2692 19468 2694
rect 19706 4700 19708 4720
rect 19708 4700 19760 4720
rect 19760 4700 19762 4720
rect 19706 4664 19762 4700
rect 20258 3712 20314 3768
rect 20074 3032 20130 3088
rect 20626 4664 20682 4720
rect 20718 4140 20774 4176
rect 20718 4120 20720 4140
rect 20720 4120 20772 4140
rect 20772 4120 20774 4140
rect 20442 2896 20498 2952
rect 22098 15272 22154 15328
rect 22190 14864 22246 14920
rect 22006 11736 22062 11792
rect 22006 9560 22062 9616
rect 23726 28314 23782 28316
rect 23806 28314 23862 28316
rect 23886 28314 23942 28316
rect 23966 28314 24022 28316
rect 23726 28262 23752 28314
rect 23752 28262 23782 28314
rect 23806 28262 23816 28314
rect 23816 28262 23862 28314
rect 23886 28262 23932 28314
rect 23932 28262 23942 28314
rect 23966 28262 23996 28314
rect 23996 28262 24022 28314
rect 23726 28260 23782 28262
rect 23806 28260 23862 28262
rect 23886 28260 23942 28262
rect 23966 28260 24022 28262
rect 23726 27226 23782 27228
rect 23806 27226 23862 27228
rect 23886 27226 23942 27228
rect 23966 27226 24022 27228
rect 23726 27174 23752 27226
rect 23752 27174 23782 27226
rect 23806 27174 23816 27226
rect 23816 27174 23862 27226
rect 23886 27174 23932 27226
rect 23932 27174 23942 27226
rect 23966 27174 23996 27226
rect 23996 27174 24022 27226
rect 23726 27172 23782 27174
rect 23806 27172 23862 27174
rect 23886 27172 23942 27174
rect 23966 27172 24022 27174
rect 23726 26138 23782 26140
rect 23806 26138 23862 26140
rect 23886 26138 23942 26140
rect 23966 26138 24022 26140
rect 23726 26086 23752 26138
rect 23752 26086 23782 26138
rect 23806 26086 23816 26138
rect 23816 26086 23862 26138
rect 23886 26086 23932 26138
rect 23932 26086 23942 26138
rect 23966 26086 23996 26138
rect 23996 26086 24022 26138
rect 23726 26084 23782 26086
rect 23806 26084 23862 26086
rect 23886 26084 23942 26086
rect 23966 26084 24022 26086
rect 23726 25050 23782 25052
rect 23806 25050 23862 25052
rect 23886 25050 23942 25052
rect 23966 25050 24022 25052
rect 23726 24998 23752 25050
rect 23752 24998 23782 25050
rect 23806 24998 23816 25050
rect 23816 24998 23862 25050
rect 23886 24998 23932 25050
rect 23932 24998 23942 25050
rect 23966 24998 23996 25050
rect 23996 24998 24022 25050
rect 23726 24996 23782 24998
rect 23806 24996 23862 24998
rect 23886 24996 23942 24998
rect 23966 24996 24022 24998
rect 23726 23962 23782 23964
rect 23806 23962 23862 23964
rect 23886 23962 23942 23964
rect 23966 23962 24022 23964
rect 23726 23910 23752 23962
rect 23752 23910 23782 23962
rect 23806 23910 23816 23962
rect 23816 23910 23862 23962
rect 23886 23910 23932 23962
rect 23932 23910 23942 23962
rect 23966 23910 23996 23962
rect 23996 23910 24022 23962
rect 23726 23908 23782 23910
rect 23806 23908 23862 23910
rect 23886 23908 23942 23910
rect 23966 23908 24022 23910
rect 23726 22874 23782 22876
rect 23806 22874 23862 22876
rect 23886 22874 23942 22876
rect 23966 22874 24022 22876
rect 23726 22822 23752 22874
rect 23752 22822 23782 22874
rect 23806 22822 23816 22874
rect 23816 22822 23862 22874
rect 23886 22822 23932 22874
rect 23932 22822 23942 22874
rect 23966 22822 23996 22874
rect 23996 22822 24022 22874
rect 23726 22820 23782 22822
rect 23806 22820 23862 22822
rect 23886 22820 23942 22822
rect 23966 22820 24022 22822
rect 23726 21786 23782 21788
rect 23806 21786 23862 21788
rect 23886 21786 23942 21788
rect 23966 21786 24022 21788
rect 23726 21734 23752 21786
rect 23752 21734 23782 21786
rect 23806 21734 23816 21786
rect 23816 21734 23862 21786
rect 23886 21734 23932 21786
rect 23932 21734 23942 21786
rect 23966 21734 23996 21786
rect 23996 21734 24022 21786
rect 23726 21732 23782 21734
rect 23806 21732 23862 21734
rect 23886 21732 23942 21734
rect 23966 21732 24022 21734
rect 23726 20698 23782 20700
rect 23806 20698 23862 20700
rect 23886 20698 23942 20700
rect 23966 20698 24022 20700
rect 23726 20646 23752 20698
rect 23752 20646 23782 20698
rect 23806 20646 23816 20698
rect 23816 20646 23862 20698
rect 23886 20646 23932 20698
rect 23932 20646 23942 20698
rect 23966 20646 23996 20698
rect 23996 20646 24022 20698
rect 23726 20644 23782 20646
rect 23806 20644 23862 20646
rect 23886 20644 23942 20646
rect 23966 20644 24022 20646
rect 22742 17060 22798 17096
rect 22742 17040 22744 17060
rect 22744 17040 22796 17060
rect 22796 17040 22798 17060
rect 23726 19610 23782 19612
rect 23806 19610 23862 19612
rect 23886 19610 23942 19612
rect 23966 19610 24022 19612
rect 23726 19558 23752 19610
rect 23752 19558 23782 19610
rect 23806 19558 23816 19610
rect 23816 19558 23862 19610
rect 23886 19558 23932 19610
rect 23932 19558 23942 19610
rect 23966 19558 23996 19610
rect 23996 19558 24022 19610
rect 23726 19556 23782 19558
rect 23806 19556 23862 19558
rect 23886 19556 23942 19558
rect 23966 19556 24022 19558
rect 23726 18522 23782 18524
rect 23806 18522 23862 18524
rect 23886 18522 23942 18524
rect 23966 18522 24022 18524
rect 23726 18470 23752 18522
rect 23752 18470 23782 18522
rect 23806 18470 23816 18522
rect 23816 18470 23862 18522
rect 23886 18470 23932 18522
rect 23932 18470 23942 18522
rect 23966 18470 23996 18522
rect 23996 18470 24022 18522
rect 23726 18468 23782 18470
rect 23806 18468 23862 18470
rect 23886 18468 23942 18470
rect 23966 18468 24022 18470
rect 23726 17434 23782 17436
rect 23806 17434 23862 17436
rect 23886 17434 23942 17436
rect 23966 17434 24022 17436
rect 23726 17382 23752 17434
rect 23752 17382 23782 17434
rect 23806 17382 23816 17434
rect 23816 17382 23862 17434
rect 23886 17382 23932 17434
rect 23932 17382 23942 17434
rect 23966 17382 23996 17434
rect 23996 17382 24022 17434
rect 23726 17380 23782 17382
rect 23806 17380 23862 17382
rect 23886 17380 23942 17382
rect 23966 17380 24022 17382
rect 23726 16346 23782 16348
rect 23806 16346 23862 16348
rect 23886 16346 23942 16348
rect 23966 16346 24022 16348
rect 23726 16294 23752 16346
rect 23752 16294 23782 16346
rect 23806 16294 23816 16346
rect 23816 16294 23862 16346
rect 23886 16294 23932 16346
rect 23932 16294 23942 16346
rect 23966 16294 23996 16346
rect 23996 16294 24022 16346
rect 23726 16292 23782 16294
rect 23806 16292 23862 16294
rect 23886 16292 23942 16294
rect 23966 16292 24022 16294
rect 23726 15258 23782 15260
rect 23806 15258 23862 15260
rect 23886 15258 23942 15260
rect 23966 15258 24022 15260
rect 23726 15206 23752 15258
rect 23752 15206 23782 15258
rect 23806 15206 23816 15258
rect 23816 15206 23862 15258
rect 23886 15206 23932 15258
rect 23932 15206 23942 15258
rect 23966 15206 23996 15258
rect 23996 15206 24022 15258
rect 23726 15204 23782 15206
rect 23806 15204 23862 15206
rect 23886 15204 23942 15206
rect 23966 15204 24022 15206
rect 24214 14900 24216 14920
rect 24216 14900 24268 14920
rect 24268 14900 24270 14920
rect 24214 14864 24270 14900
rect 23726 14170 23782 14172
rect 23806 14170 23862 14172
rect 23886 14170 23942 14172
rect 23966 14170 24022 14172
rect 23726 14118 23752 14170
rect 23752 14118 23782 14170
rect 23806 14118 23816 14170
rect 23816 14118 23862 14170
rect 23886 14118 23932 14170
rect 23932 14118 23942 14170
rect 23966 14118 23996 14170
rect 23996 14118 24022 14170
rect 23726 14116 23782 14118
rect 23806 14116 23862 14118
rect 23886 14116 23942 14118
rect 23966 14116 24022 14118
rect 23726 13082 23782 13084
rect 23806 13082 23862 13084
rect 23886 13082 23942 13084
rect 23966 13082 24022 13084
rect 23726 13030 23752 13082
rect 23752 13030 23782 13082
rect 23806 13030 23816 13082
rect 23816 13030 23862 13082
rect 23886 13030 23932 13082
rect 23932 13030 23942 13082
rect 23966 13030 23996 13082
rect 23996 13030 24022 13082
rect 23726 13028 23782 13030
rect 23806 13028 23862 13030
rect 23886 13028 23942 13030
rect 23966 13028 24022 13030
rect 23202 11192 23258 11248
rect 23018 7948 23074 7984
rect 23018 7928 23020 7948
rect 23020 7928 23072 7948
rect 23072 7928 23074 7948
rect 22834 7792 22890 7848
rect 23726 11994 23782 11996
rect 23806 11994 23862 11996
rect 23886 11994 23942 11996
rect 23966 11994 24022 11996
rect 23726 11942 23752 11994
rect 23752 11942 23782 11994
rect 23806 11942 23816 11994
rect 23816 11942 23862 11994
rect 23886 11942 23932 11994
rect 23932 11942 23942 11994
rect 23966 11942 23996 11994
rect 23996 11942 24022 11994
rect 23726 11940 23782 11942
rect 23806 11940 23862 11942
rect 23886 11940 23942 11942
rect 23966 11940 24022 11942
rect 23754 11212 23810 11248
rect 24214 11736 24270 11792
rect 23754 11192 23756 11212
rect 23756 11192 23808 11212
rect 23808 11192 23810 11212
rect 23726 10906 23782 10908
rect 23806 10906 23862 10908
rect 23886 10906 23942 10908
rect 23966 10906 24022 10908
rect 23726 10854 23752 10906
rect 23752 10854 23782 10906
rect 23806 10854 23816 10906
rect 23816 10854 23862 10906
rect 23886 10854 23932 10906
rect 23932 10854 23942 10906
rect 23966 10854 23996 10906
rect 23996 10854 24022 10906
rect 23726 10852 23782 10854
rect 23806 10852 23862 10854
rect 23886 10852 23942 10854
rect 23966 10852 24022 10854
rect 23726 9818 23782 9820
rect 23806 9818 23862 9820
rect 23886 9818 23942 9820
rect 23966 9818 24022 9820
rect 23726 9766 23752 9818
rect 23752 9766 23782 9818
rect 23806 9766 23816 9818
rect 23816 9766 23862 9818
rect 23886 9766 23932 9818
rect 23932 9766 23942 9818
rect 23966 9766 23996 9818
rect 23996 9766 24022 9818
rect 23726 9764 23782 9766
rect 23806 9764 23862 9766
rect 23886 9764 23942 9766
rect 23966 9764 24022 9766
rect 23726 8730 23782 8732
rect 23806 8730 23862 8732
rect 23886 8730 23942 8732
rect 23966 8730 24022 8732
rect 23726 8678 23752 8730
rect 23752 8678 23782 8730
rect 23806 8678 23816 8730
rect 23816 8678 23862 8730
rect 23886 8678 23932 8730
rect 23932 8678 23942 8730
rect 23966 8678 23996 8730
rect 23996 8678 24022 8730
rect 23726 8676 23782 8678
rect 23806 8676 23862 8678
rect 23886 8676 23942 8678
rect 23966 8676 24022 8678
rect 23726 7642 23782 7644
rect 23806 7642 23862 7644
rect 23886 7642 23942 7644
rect 23966 7642 24022 7644
rect 23726 7590 23752 7642
rect 23752 7590 23782 7642
rect 23806 7590 23816 7642
rect 23816 7590 23862 7642
rect 23886 7590 23932 7642
rect 23932 7590 23942 7642
rect 23966 7590 23996 7642
rect 23996 7590 24022 7642
rect 23726 7588 23782 7590
rect 23806 7588 23862 7590
rect 23886 7588 23942 7590
rect 23966 7588 24022 7590
rect 23726 6554 23782 6556
rect 23806 6554 23862 6556
rect 23886 6554 23942 6556
rect 23966 6554 24022 6556
rect 23726 6502 23752 6554
rect 23752 6502 23782 6554
rect 23806 6502 23816 6554
rect 23816 6502 23862 6554
rect 23886 6502 23932 6554
rect 23932 6502 23942 6554
rect 23966 6502 23996 6554
rect 23996 6502 24022 6554
rect 23726 6500 23782 6502
rect 23806 6500 23862 6502
rect 23886 6500 23942 6502
rect 23966 6500 24022 6502
rect 23110 6196 23112 6216
rect 23112 6196 23164 6216
rect 23164 6196 23166 6216
rect 23110 6160 23166 6196
rect 23018 4392 23074 4448
rect 23726 5466 23782 5468
rect 23806 5466 23862 5468
rect 23886 5466 23942 5468
rect 23966 5466 24022 5468
rect 23726 5414 23752 5466
rect 23752 5414 23782 5466
rect 23806 5414 23816 5466
rect 23816 5414 23862 5466
rect 23886 5414 23932 5466
rect 23932 5414 23942 5466
rect 23966 5414 23996 5466
rect 23996 5414 24022 5466
rect 23726 5412 23782 5414
rect 23806 5412 23862 5414
rect 23886 5412 23942 5414
rect 23966 5412 24022 5414
rect 23726 4378 23782 4380
rect 23806 4378 23862 4380
rect 23886 4378 23942 4380
rect 23966 4378 24022 4380
rect 23726 4326 23752 4378
rect 23752 4326 23782 4378
rect 23806 4326 23816 4378
rect 23816 4326 23862 4378
rect 23886 4326 23932 4378
rect 23932 4326 23942 4378
rect 23966 4326 23996 4378
rect 23996 4326 24022 4378
rect 23726 4324 23782 4326
rect 23806 4324 23862 4326
rect 23886 4324 23942 4326
rect 23966 4324 24022 4326
rect 23938 4004 23994 4040
rect 23938 3984 23940 4004
rect 23940 3984 23992 4004
rect 23992 3984 23994 4004
rect 24398 3712 24454 3768
rect 23726 3290 23782 3292
rect 23806 3290 23862 3292
rect 23886 3290 23942 3292
rect 23966 3290 24022 3292
rect 23726 3238 23752 3290
rect 23752 3238 23782 3290
rect 23806 3238 23816 3290
rect 23816 3238 23862 3290
rect 23886 3238 23932 3290
rect 23932 3238 23942 3290
rect 23966 3238 23996 3290
rect 23996 3238 24022 3290
rect 23726 3236 23782 3238
rect 23806 3236 23862 3238
rect 23886 3236 23942 3238
rect 23966 3236 24022 3238
rect 23726 2202 23782 2204
rect 23806 2202 23862 2204
rect 23886 2202 23942 2204
rect 23966 2202 24022 2204
rect 23726 2150 23752 2202
rect 23752 2150 23782 2202
rect 23806 2150 23816 2202
rect 23816 2150 23862 2202
rect 23886 2150 23932 2202
rect 23932 2150 23942 2202
rect 23966 2150 23996 2202
rect 23996 2150 24022 2202
rect 23726 2148 23782 2150
rect 23806 2148 23862 2150
rect 23886 2148 23942 2150
rect 23966 2148 24022 2150
rect 24858 20440 24914 20496
rect 24950 17040 25006 17096
rect 25134 22480 25190 22536
rect 26146 30640 26202 30696
rect 26054 29280 26110 29336
rect 25686 19352 25742 19408
rect 25502 17740 25558 17776
rect 25502 17720 25504 17740
rect 25504 17720 25556 17740
rect 25556 17720 25558 17740
rect 25134 15680 25190 15736
rect 25594 15680 25650 15736
rect 24766 6160 24822 6216
rect 26146 27920 26202 27976
rect 26330 23432 26386 23488
rect 26146 17040 26202 17096
rect 26146 14320 26202 14376
rect 26146 6840 26202 6896
rect 25962 1400 26018 1456
rect 26882 28600 26938 28656
rect 26882 25900 26938 25936
rect 26882 25880 26884 25900
rect 26884 25880 26936 25900
rect 26936 25880 26938 25900
rect 26790 23840 26846 23896
rect 26606 23604 26608 23624
rect 26608 23604 26660 23624
rect 26660 23604 26662 23624
rect 26606 23568 26662 23604
rect 26974 25200 27030 25256
rect 26974 23160 27030 23216
rect 26882 18400 26938 18456
rect 26882 15000 26938 15056
rect 26882 11600 26938 11656
rect 26146 3984 26202 4040
rect 26790 10240 26846 10296
rect 26698 9560 26754 9616
rect 26698 7520 26754 7576
rect 27710 26560 27766 26616
rect 26790 4120 26846 4176
rect 26882 3440 26938 3496
rect 26514 2080 26570 2136
rect 27618 21936 27674 21992
rect 27526 21120 27582 21176
rect 27526 19760 27582 19816
rect 27526 8880 27582 8936
rect 27802 12960 27858 13016
rect 27710 12300 27766 12336
rect 27710 12280 27712 12300
rect 27712 12280 27764 12300
rect 27764 12280 27766 12300
rect 27710 8900 27766 8936
rect 27710 8880 27712 8900
rect 27712 8880 27764 8900
rect 27764 8880 27766 8900
rect 27710 6160 27766 6216
rect 27526 4800 27582 4856
rect 26054 720 26110 776
<< metal3 >>
rect 0 30698 800 30728
rect 2865 30698 2931 30701
rect 0 30696 2931 30698
rect 0 30640 2870 30696
rect 2926 30640 2931 30696
rect 0 30638 2931 30640
rect 0 30608 800 30638
rect 2865 30635 2931 30638
rect 26141 30698 26207 30701
rect 28780 30698 29580 30728
rect 26141 30696 29580 30698
rect 26141 30640 26146 30696
rect 26202 30640 29580 30696
rect 26141 30638 29580 30640
rect 26141 30635 26207 30638
rect 28780 30608 29580 30638
rect 5498 29408 5818 29409
rect 0 29338 800 29368
rect 5498 29344 5506 29408
rect 5570 29344 5586 29408
rect 5650 29344 5666 29408
rect 5730 29344 5746 29408
rect 5810 29344 5818 29408
rect 5498 29343 5818 29344
rect 14606 29408 14926 29409
rect 14606 29344 14614 29408
rect 14678 29344 14694 29408
rect 14758 29344 14774 29408
rect 14838 29344 14854 29408
rect 14918 29344 14926 29408
rect 14606 29343 14926 29344
rect 23714 29408 24034 29409
rect 23714 29344 23722 29408
rect 23786 29344 23802 29408
rect 23866 29344 23882 29408
rect 23946 29344 23962 29408
rect 24026 29344 24034 29408
rect 23714 29343 24034 29344
rect 1853 29338 1919 29341
rect 0 29336 1919 29338
rect 0 29280 1858 29336
rect 1914 29280 1919 29336
rect 0 29278 1919 29280
rect 0 29248 800 29278
rect 1853 29275 1919 29278
rect 26049 29338 26115 29341
rect 28780 29338 29580 29368
rect 26049 29336 29580 29338
rect 26049 29280 26054 29336
rect 26110 29280 29580 29336
rect 26049 29278 29580 29280
rect 26049 29275 26115 29278
rect 28780 29248 29580 29278
rect 10052 28864 10372 28865
rect 10052 28800 10060 28864
rect 10124 28800 10140 28864
rect 10204 28800 10220 28864
rect 10284 28800 10300 28864
rect 10364 28800 10372 28864
rect 10052 28799 10372 28800
rect 19160 28864 19480 28865
rect 19160 28800 19168 28864
rect 19232 28800 19248 28864
rect 19312 28800 19328 28864
rect 19392 28800 19408 28864
rect 19472 28800 19480 28864
rect 19160 28799 19480 28800
rect 0 28658 800 28688
rect 2129 28658 2195 28661
rect 0 28656 2195 28658
rect 0 28600 2134 28656
rect 2190 28600 2195 28656
rect 0 28598 2195 28600
rect 0 28568 800 28598
rect 2129 28595 2195 28598
rect 7465 28658 7531 28661
rect 8569 28658 8635 28661
rect 9857 28660 9923 28661
rect 9806 28658 9812 28660
rect 7465 28656 8635 28658
rect 7465 28600 7470 28656
rect 7526 28600 8574 28656
rect 8630 28600 8635 28656
rect 7465 28598 8635 28600
rect 9766 28598 9812 28658
rect 9876 28656 9923 28660
rect 9918 28600 9923 28656
rect 7465 28595 7531 28598
rect 8569 28595 8635 28598
rect 9806 28596 9812 28598
rect 9876 28596 9923 28600
rect 9857 28595 9923 28596
rect 26877 28658 26943 28661
rect 28780 28658 29580 28688
rect 26877 28656 29580 28658
rect 26877 28600 26882 28656
rect 26938 28600 29580 28656
rect 26877 28598 29580 28600
rect 26877 28595 26943 28598
rect 28780 28568 29580 28598
rect 5498 28320 5818 28321
rect 5498 28256 5506 28320
rect 5570 28256 5586 28320
rect 5650 28256 5666 28320
rect 5730 28256 5746 28320
rect 5810 28256 5818 28320
rect 5498 28255 5818 28256
rect 14606 28320 14926 28321
rect 14606 28256 14614 28320
rect 14678 28256 14694 28320
rect 14758 28256 14774 28320
rect 14838 28256 14854 28320
rect 14918 28256 14926 28320
rect 14606 28255 14926 28256
rect 23714 28320 24034 28321
rect 23714 28256 23722 28320
rect 23786 28256 23802 28320
rect 23866 28256 23882 28320
rect 23946 28256 23962 28320
rect 24026 28256 24034 28320
rect 23714 28255 24034 28256
rect 0 27978 800 28008
rect 1393 27978 1459 27981
rect 0 27976 1459 27978
rect 0 27920 1398 27976
rect 1454 27920 1459 27976
rect 0 27918 1459 27920
rect 0 27888 800 27918
rect 1393 27915 1459 27918
rect 26141 27978 26207 27981
rect 28780 27978 29580 28008
rect 26141 27976 29580 27978
rect 26141 27920 26146 27976
rect 26202 27920 29580 27976
rect 26141 27918 29580 27920
rect 26141 27915 26207 27918
rect 28780 27888 29580 27918
rect 10052 27776 10372 27777
rect 10052 27712 10060 27776
rect 10124 27712 10140 27776
rect 10204 27712 10220 27776
rect 10284 27712 10300 27776
rect 10364 27712 10372 27776
rect 10052 27711 10372 27712
rect 19160 27776 19480 27777
rect 19160 27712 19168 27776
rect 19232 27712 19248 27776
rect 19312 27712 19328 27776
rect 19392 27712 19408 27776
rect 19472 27712 19480 27776
rect 19160 27711 19480 27712
rect 10501 27570 10567 27573
rect 15101 27570 15167 27573
rect 10501 27568 15167 27570
rect 10501 27512 10506 27568
rect 10562 27512 15106 27568
rect 15162 27512 15167 27568
rect 10501 27510 15167 27512
rect 10501 27507 10567 27510
rect 15101 27507 15167 27510
rect 5498 27232 5818 27233
rect 5498 27168 5506 27232
rect 5570 27168 5586 27232
rect 5650 27168 5666 27232
rect 5730 27168 5746 27232
rect 5810 27168 5818 27232
rect 5498 27167 5818 27168
rect 14606 27232 14926 27233
rect 14606 27168 14614 27232
rect 14678 27168 14694 27232
rect 14758 27168 14774 27232
rect 14838 27168 14854 27232
rect 14918 27168 14926 27232
rect 14606 27167 14926 27168
rect 23714 27232 24034 27233
rect 23714 27168 23722 27232
rect 23786 27168 23802 27232
rect 23866 27168 23882 27232
rect 23946 27168 23962 27232
rect 24026 27168 24034 27232
rect 23714 27167 24034 27168
rect 9765 27162 9831 27165
rect 9630 27160 9831 27162
rect 9630 27104 9770 27160
rect 9826 27104 9831 27160
rect 9630 27102 9831 27104
rect 9630 26893 9690 27102
rect 9765 27099 9831 27102
rect 9630 26888 9739 26893
rect 9630 26832 9678 26888
rect 9734 26832 9739 26888
rect 9630 26830 9739 26832
rect 9673 26827 9739 26830
rect 10052 26688 10372 26689
rect 0 26618 800 26648
rect 10052 26624 10060 26688
rect 10124 26624 10140 26688
rect 10204 26624 10220 26688
rect 10284 26624 10300 26688
rect 10364 26624 10372 26688
rect 10052 26623 10372 26624
rect 19160 26688 19480 26689
rect 19160 26624 19168 26688
rect 19232 26624 19248 26688
rect 19312 26624 19328 26688
rect 19392 26624 19408 26688
rect 19472 26624 19480 26688
rect 19160 26623 19480 26624
rect 1945 26618 2011 26621
rect 0 26616 2011 26618
rect 0 26560 1950 26616
rect 2006 26560 2011 26616
rect 0 26558 2011 26560
rect 0 26528 800 26558
rect 1945 26555 2011 26558
rect 27705 26618 27771 26621
rect 28780 26618 29580 26648
rect 27705 26616 29580 26618
rect 27705 26560 27710 26616
rect 27766 26560 29580 26616
rect 27705 26558 29580 26560
rect 27705 26555 27771 26558
rect 28780 26528 29580 26558
rect 5498 26144 5818 26145
rect 5498 26080 5506 26144
rect 5570 26080 5586 26144
rect 5650 26080 5666 26144
rect 5730 26080 5746 26144
rect 5810 26080 5818 26144
rect 5498 26079 5818 26080
rect 14606 26144 14926 26145
rect 14606 26080 14614 26144
rect 14678 26080 14694 26144
rect 14758 26080 14774 26144
rect 14838 26080 14854 26144
rect 14918 26080 14926 26144
rect 14606 26079 14926 26080
rect 23714 26144 24034 26145
rect 23714 26080 23722 26144
rect 23786 26080 23802 26144
rect 23866 26080 23882 26144
rect 23946 26080 23962 26144
rect 24026 26080 24034 26144
rect 23714 26079 24034 26080
rect 0 25938 800 25968
rect 1669 25938 1735 25941
rect 0 25936 1735 25938
rect 0 25880 1674 25936
rect 1730 25880 1735 25936
rect 0 25878 1735 25880
rect 0 25848 800 25878
rect 1669 25875 1735 25878
rect 26877 25938 26943 25941
rect 28780 25938 29580 25968
rect 26877 25936 29580 25938
rect 26877 25880 26882 25936
rect 26938 25880 29580 25936
rect 26877 25878 29580 25880
rect 26877 25875 26943 25878
rect 28780 25848 29580 25878
rect 10052 25600 10372 25601
rect 10052 25536 10060 25600
rect 10124 25536 10140 25600
rect 10204 25536 10220 25600
rect 10284 25536 10300 25600
rect 10364 25536 10372 25600
rect 10052 25535 10372 25536
rect 19160 25600 19480 25601
rect 19160 25536 19168 25600
rect 19232 25536 19248 25600
rect 19312 25536 19328 25600
rect 19392 25536 19408 25600
rect 19472 25536 19480 25600
rect 19160 25535 19480 25536
rect 10961 25394 11027 25397
rect 13445 25394 13511 25397
rect 10961 25392 13511 25394
rect 10961 25336 10966 25392
rect 11022 25336 13450 25392
rect 13506 25336 13511 25392
rect 10961 25334 13511 25336
rect 10961 25331 11027 25334
rect 13445 25331 13511 25334
rect 0 25258 800 25288
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25168 800 25198
rect 1393 25195 1459 25198
rect 26969 25258 27035 25261
rect 28780 25258 29580 25288
rect 26969 25256 29580 25258
rect 26969 25200 26974 25256
rect 27030 25200 29580 25256
rect 26969 25198 29580 25200
rect 26969 25195 27035 25198
rect 28780 25168 29580 25198
rect 5498 25056 5818 25057
rect 5498 24992 5506 25056
rect 5570 24992 5586 25056
rect 5650 24992 5666 25056
rect 5730 24992 5746 25056
rect 5810 24992 5818 25056
rect 5498 24991 5818 24992
rect 14606 25056 14926 25057
rect 14606 24992 14614 25056
rect 14678 24992 14694 25056
rect 14758 24992 14774 25056
rect 14838 24992 14854 25056
rect 14918 24992 14926 25056
rect 14606 24991 14926 24992
rect 23714 25056 24034 25057
rect 23714 24992 23722 25056
rect 23786 24992 23802 25056
rect 23866 24992 23882 25056
rect 23946 24992 23962 25056
rect 24026 24992 24034 25056
rect 23714 24991 24034 24992
rect 14273 24850 14339 24853
rect 14917 24850 14983 24853
rect 15929 24850 15995 24853
rect 14273 24848 15995 24850
rect 14273 24792 14278 24848
rect 14334 24792 14922 24848
rect 14978 24792 15934 24848
rect 15990 24792 15995 24848
rect 14273 24790 15995 24792
rect 14273 24787 14339 24790
rect 14917 24787 14983 24790
rect 15929 24787 15995 24790
rect 12341 24714 12407 24717
rect 15653 24714 15719 24717
rect 12341 24712 15719 24714
rect 12341 24656 12346 24712
rect 12402 24656 15658 24712
rect 15714 24656 15719 24712
rect 12341 24654 15719 24656
rect 12341 24651 12407 24654
rect 15653 24651 15719 24654
rect 10052 24512 10372 24513
rect 10052 24448 10060 24512
rect 10124 24448 10140 24512
rect 10204 24448 10220 24512
rect 10284 24448 10300 24512
rect 10364 24448 10372 24512
rect 10052 24447 10372 24448
rect 19160 24512 19480 24513
rect 19160 24448 19168 24512
rect 19232 24448 19248 24512
rect 19312 24448 19328 24512
rect 19392 24448 19408 24512
rect 19472 24448 19480 24512
rect 19160 24447 19480 24448
rect 9857 24172 9923 24173
rect 9806 24108 9812 24172
rect 9876 24170 9923 24172
rect 9876 24168 9968 24170
rect 9918 24112 9968 24168
rect 9876 24110 9968 24112
rect 9876 24108 9923 24110
rect 9857 24107 9923 24108
rect 5498 23968 5818 23969
rect 0 23898 800 23928
rect 5498 23904 5506 23968
rect 5570 23904 5586 23968
rect 5650 23904 5666 23968
rect 5730 23904 5746 23968
rect 5810 23904 5818 23968
rect 5498 23903 5818 23904
rect 14606 23968 14926 23969
rect 14606 23904 14614 23968
rect 14678 23904 14694 23968
rect 14758 23904 14774 23968
rect 14838 23904 14854 23968
rect 14918 23904 14926 23968
rect 14606 23903 14926 23904
rect 23714 23968 24034 23969
rect 23714 23904 23722 23968
rect 23786 23904 23802 23968
rect 23866 23904 23882 23968
rect 23946 23904 23962 23968
rect 24026 23904 24034 23968
rect 23714 23903 24034 23904
rect 1669 23898 1735 23901
rect 0 23896 1735 23898
rect 0 23840 1674 23896
rect 1730 23840 1735 23896
rect 0 23838 1735 23840
rect 0 23808 800 23838
rect 1669 23835 1735 23838
rect 26785 23898 26851 23901
rect 28780 23898 29580 23928
rect 26785 23896 29580 23898
rect 26785 23840 26790 23896
rect 26846 23840 29580 23896
rect 26785 23838 29580 23840
rect 26785 23835 26851 23838
rect 28780 23808 29580 23838
rect 21265 23626 21331 23629
rect 26601 23626 26667 23629
rect 21265 23624 26667 23626
rect 21265 23568 21270 23624
rect 21326 23568 26606 23624
rect 26662 23568 26667 23624
rect 21265 23566 26667 23568
rect 21265 23563 21331 23566
rect 26601 23563 26667 23566
rect 26325 23492 26391 23493
rect 26325 23488 26372 23492
rect 26436 23490 26442 23492
rect 26325 23432 26330 23488
rect 26325 23428 26372 23432
rect 26436 23430 26482 23490
rect 26436 23428 26442 23430
rect 26325 23427 26391 23428
rect 10052 23424 10372 23425
rect 10052 23360 10060 23424
rect 10124 23360 10140 23424
rect 10204 23360 10220 23424
rect 10284 23360 10300 23424
rect 10364 23360 10372 23424
rect 10052 23359 10372 23360
rect 19160 23424 19480 23425
rect 19160 23360 19168 23424
rect 19232 23360 19248 23424
rect 19312 23360 19328 23424
rect 19392 23360 19408 23424
rect 19472 23360 19480 23424
rect 19160 23359 19480 23360
rect 14457 23354 14523 23357
rect 18781 23354 18847 23357
rect 14457 23352 18847 23354
rect 14457 23296 14462 23352
rect 14518 23296 18786 23352
rect 18842 23296 18847 23352
rect 14457 23294 18847 23296
rect 14457 23291 14523 23294
rect 18781 23291 18847 23294
rect 0 23218 800 23248
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23128 800 23158
rect 1853 23155 1919 23158
rect 10685 23218 10751 23221
rect 18689 23218 18755 23221
rect 10685 23216 18755 23218
rect 10685 23160 10690 23216
rect 10746 23160 18694 23216
rect 18750 23160 18755 23216
rect 10685 23158 18755 23160
rect 10685 23155 10751 23158
rect 18689 23155 18755 23158
rect 26969 23218 27035 23221
rect 28780 23218 29580 23248
rect 26969 23216 29580 23218
rect 26969 23160 26974 23216
rect 27030 23160 29580 23216
rect 26969 23158 29580 23160
rect 26969 23155 27035 23158
rect 28780 23128 29580 23158
rect 14825 23082 14891 23085
rect 19149 23082 19215 23085
rect 14825 23080 19215 23082
rect 14825 23024 14830 23080
rect 14886 23024 19154 23080
rect 19210 23024 19215 23080
rect 14825 23022 19215 23024
rect 14825 23019 14891 23022
rect 19149 23019 19215 23022
rect 5498 22880 5818 22881
rect 5498 22816 5506 22880
rect 5570 22816 5586 22880
rect 5650 22816 5666 22880
rect 5730 22816 5746 22880
rect 5810 22816 5818 22880
rect 5498 22815 5818 22816
rect 14606 22880 14926 22881
rect 14606 22816 14614 22880
rect 14678 22816 14694 22880
rect 14758 22816 14774 22880
rect 14838 22816 14854 22880
rect 14918 22816 14926 22880
rect 14606 22815 14926 22816
rect 23714 22880 24034 22881
rect 23714 22816 23722 22880
rect 23786 22816 23802 22880
rect 23866 22816 23882 22880
rect 23946 22816 23962 22880
rect 24026 22816 24034 22880
rect 23714 22815 24034 22816
rect 0 22538 800 22568
rect 2037 22538 2103 22541
rect 0 22536 2103 22538
rect 0 22480 2042 22536
rect 2098 22480 2103 22536
rect 0 22478 2103 22480
rect 0 22448 800 22478
rect 2037 22475 2103 22478
rect 25129 22538 25195 22541
rect 28780 22538 29580 22568
rect 25129 22536 29580 22538
rect 25129 22480 25134 22536
rect 25190 22480 29580 22536
rect 25129 22478 29580 22480
rect 25129 22475 25195 22478
rect 28780 22448 29580 22478
rect 10052 22336 10372 22337
rect 10052 22272 10060 22336
rect 10124 22272 10140 22336
rect 10204 22272 10220 22336
rect 10284 22272 10300 22336
rect 10364 22272 10372 22336
rect 10052 22271 10372 22272
rect 19160 22336 19480 22337
rect 19160 22272 19168 22336
rect 19232 22272 19248 22336
rect 19312 22272 19328 22336
rect 19392 22272 19408 22336
rect 19472 22272 19480 22336
rect 19160 22271 19480 22272
rect 18229 22130 18295 22133
rect 20897 22130 20963 22133
rect 18229 22128 20963 22130
rect 18229 22072 18234 22128
rect 18290 22072 20902 22128
rect 20958 22072 20963 22128
rect 18229 22070 20963 22072
rect 18229 22067 18295 22070
rect 20897 22067 20963 22070
rect 13261 21994 13327 21997
rect 27613 21994 27679 21997
rect 13261 21992 27679 21994
rect 13261 21936 13266 21992
rect 13322 21936 27618 21992
rect 27674 21936 27679 21992
rect 13261 21934 27679 21936
rect 13261 21931 13327 21934
rect 27613 21931 27679 21934
rect 5498 21792 5818 21793
rect 5498 21728 5506 21792
rect 5570 21728 5586 21792
rect 5650 21728 5666 21792
rect 5730 21728 5746 21792
rect 5810 21728 5818 21792
rect 5498 21727 5818 21728
rect 14606 21792 14926 21793
rect 14606 21728 14614 21792
rect 14678 21728 14694 21792
rect 14758 21728 14774 21792
rect 14838 21728 14854 21792
rect 14918 21728 14926 21792
rect 14606 21727 14926 21728
rect 23714 21792 24034 21793
rect 23714 21728 23722 21792
rect 23786 21728 23802 21792
rect 23866 21728 23882 21792
rect 23946 21728 23962 21792
rect 24026 21728 24034 21792
rect 23714 21727 24034 21728
rect 9673 21586 9739 21589
rect 18229 21586 18295 21589
rect 9673 21584 18295 21586
rect 9673 21528 9678 21584
rect 9734 21528 18234 21584
rect 18290 21528 18295 21584
rect 9673 21526 18295 21528
rect 9673 21523 9739 21526
rect 18229 21523 18295 21526
rect 18229 21450 18295 21453
rect 19241 21450 19307 21453
rect 18229 21448 19307 21450
rect 18229 21392 18234 21448
rect 18290 21392 19246 21448
rect 19302 21392 19307 21448
rect 18229 21390 19307 21392
rect 18229 21387 18295 21390
rect 19241 21387 19307 21390
rect 4245 21314 4311 21317
rect 5441 21314 5507 21317
rect 6913 21314 6979 21317
rect 4245 21312 6979 21314
rect 4245 21256 4250 21312
rect 4306 21256 5446 21312
rect 5502 21256 6918 21312
rect 6974 21256 6979 21312
rect 4245 21254 6979 21256
rect 4245 21251 4311 21254
rect 5441 21251 5507 21254
rect 6913 21251 6979 21254
rect 13261 21314 13327 21317
rect 14089 21314 14155 21317
rect 13261 21312 14155 21314
rect 13261 21256 13266 21312
rect 13322 21256 14094 21312
rect 14150 21256 14155 21312
rect 13261 21254 14155 21256
rect 13261 21251 13327 21254
rect 14089 21251 14155 21254
rect 10052 21248 10372 21249
rect 0 21178 800 21208
rect 10052 21184 10060 21248
rect 10124 21184 10140 21248
rect 10204 21184 10220 21248
rect 10284 21184 10300 21248
rect 10364 21184 10372 21248
rect 10052 21183 10372 21184
rect 19160 21248 19480 21249
rect 19160 21184 19168 21248
rect 19232 21184 19248 21248
rect 19312 21184 19328 21248
rect 19392 21184 19408 21248
rect 19472 21184 19480 21248
rect 19160 21183 19480 21184
rect 1945 21178 2011 21181
rect 0 21176 2011 21178
rect 0 21120 1950 21176
rect 2006 21120 2011 21176
rect 0 21118 2011 21120
rect 0 21088 800 21118
rect 1945 21115 2011 21118
rect 27521 21178 27587 21181
rect 28780 21178 29580 21208
rect 27521 21176 29580 21178
rect 27521 21120 27526 21176
rect 27582 21120 29580 21176
rect 27521 21118 29580 21120
rect 27521 21115 27587 21118
rect 28780 21088 29580 21118
rect 5498 20704 5818 20705
rect 5498 20640 5506 20704
rect 5570 20640 5586 20704
rect 5650 20640 5666 20704
rect 5730 20640 5746 20704
rect 5810 20640 5818 20704
rect 5498 20639 5818 20640
rect 14606 20704 14926 20705
rect 14606 20640 14614 20704
rect 14678 20640 14694 20704
rect 14758 20640 14774 20704
rect 14838 20640 14854 20704
rect 14918 20640 14926 20704
rect 14606 20639 14926 20640
rect 23714 20704 24034 20705
rect 23714 20640 23722 20704
rect 23786 20640 23802 20704
rect 23866 20640 23882 20704
rect 23946 20640 23962 20704
rect 24026 20640 24034 20704
rect 23714 20639 24034 20640
rect 0 20498 800 20528
rect 1669 20498 1735 20501
rect 0 20496 1735 20498
rect 0 20440 1674 20496
rect 1730 20440 1735 20496
rect 0 20438 1735 20440
rect 0 20408 800 20438
rect 1669 20435 1735 20438
rect 24853 20498 24919 20501
rect 28780 20498 29580 20528
rect 24853 20496 29580 20498
rect 24853 20440 24858 20496
rect 24914 20440 29580 20496
rect 24853 20438 29580 20440
rect 24853 20435 24919 20438
rect 28780 20408 29580 20438
rect 10052 20160 10372 20161
rect 10052 20096 10060 20160
rect 10124 20096 10140 20160
rect 10204 20096 10220 20160
rect 10284 20096 10300 20160
rect 10364 20096 10372 20160
rect 10052 20095 10372 20096
rect 19160 20160 19480 20161
rect 19160 20096 19168 20160
rect 19232 20096 19248 20160
rect 19312 20096 19328 20160
rect 19392 20096 19408 20160
rect 19472 20096 19480 20160
rect 19160 20095 19480 20096
rect 5441 19954 5507 19957
rect 8477 19954 8543 19957
rect 5441 19952 8543 19954
rect 5441 19896 5446 19952
rect 5502 19896 8482 19952
rect 8538 19896 8543 19952
rect 5441 19894 8543 19896
rect 5441 19891 5507 19894
rect 8477 19891 8543 19894
rect 0 19818 800 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 800 19758
rect 1945 19755 2011 19758
rect 27521 19818 27587 19821
rect 28780 19818 29580 19848
rect 27521 19816 29580 19818
rect 27521 19760 27526 19816
rect 27582 19760 29580 19816
rect 27521 19758 29580 19760
rect 27521 19755 27587 19758
rect 28780 19728 29580 19758
rect 5498 19616 5818 19617
rect 5498 19552 5506 19616
rect 5570 19552 5586 19616
rect 5650 19552 5666 19616
rect 5730 19552 5746 19616
rect 5810 19552 5818 19616
rect 5498 19551 5818 19552
rect 14606 19616 14926 19617
rect 14606 19552 14614 19616
rect 14678 19552 14694 19616
rect 14758 19552 14774 19616
rect 14838 19552 14854 19616
rect 14918 19552 14926 19616
rect 14606 19551 14926 19552
rect 23714 19616 24034 19617
rect 23714 19552 23722 19616
rect 23786 19552 23802 19616
rect 23866 19552 23882 19616
rect 23946 19552 23962 19616
rect 24026 19552 24034 19616
rect 23714 19551 24034 19552
rect 19977 19410 20043 19413
rect 25681 19410 25747 19413
rect 19977 19408 25747 19410
rect 19977 19352 19982 19408
rect 20038 19352 25686 19408
rect 25742 19352 25747 19408
rect 19977 19350 25747 19352
rect 19977 19347 20043 19350
rect 25681 19347 25747 19350
rect 4705 19274 4771 19277
rect 7465 19274 7531 19277
rect 4705 19272 7531 19274
rect 4705 19216 4710 19272
rect 4766 19216 7470 19272
rect 7526 19216 7531 19272
rect 4705 19214 7531 19216
rect 4705 19211 4771 19214
rect 7465 19211 7531 19214
rect 9806 19212 9812 19276
rect 9876 19274 9882 19276
rect 10041 19274 10107 19277
rect 9876 19272 10107 19274
rect 9876 19216 10046 19272
rect 10102 19216 10107 19272
rect 9876 19214 10107 19216
rect 9876 19212 9882 19214
rect 10041 19211 10107 19214
rect 11881 19274 11947 19277
rect 15469 19274 15535 19277
rect 11881 19272 15535 19274
rect 11881 19216 11886 19272
rect 11942 19216 15474 19272
rect 15530 19216 15535 19272
rect 11881 19214 15535 19216
rect 11881 19211 11947 19214
rect 15469 19211 15535 19214
rect 10052 19072 10372 19073
rect 10052 19008 10060 19072
rect 10124 19008 10140 19072
rect 10204 19008 10220 19072
rect 10284 19008 10300 19072
rect 10364 19008 10372 19072
rect 10052 19007 10372 19008
rect 19160 19072 19480 19073
rect 19160 19008 19168 19072
rect 19232 19008 19248 19072
rect 19312 19008 19328 19072
rect 19392 19008 19408 19072
rect 19472 19008 19480 19072
rect 19160 19007 19480 19008
rect 12341 18866 12407 18869
rect 13169 18866 13235 18869
rect 14457 18866 14523 18869
rect 12341 18864 14523 18866
rect 12341 18808 12346 18864
rect 12402 18808 13174 18864
rect 13230 18808 14462 18864
rect 14518 18808 14523 18864
rect 12341 18806 14523 18808
rect 12341 18803 12407 18806
rect 13169 18803 13235 18806
rect 14457 18803 14523 18806
rect 14641 18866 14707 18869
rect 14641 18864 17648 18866
rect 14641 18808 14646 18864
rect 14702 18808 17648 18864
rect 14641 18806 17648 18808
rect 14641 18803 14707 18806
rect 17588 18733 17648 18806
rect 10225 18730 10291 18733
rect 15285 18730 15351 18733
rect 17125 18730 17191 18733
rect 10225 18728 17191 18730
rect 10225 18672 10230 18728
rect 10286 18672 15290 18728
rect 15346 18672 17130 18728
rect 17186 18672 17191 18728
rect 10225 18670 17191 18672
rect 10225 18667 10291 18670
rect 15285 18667 15351 18670
rect 17125 18667 17191 18670
rect 17585 18728 17651 18733
rect 17585 18672 17590 18728
rect 17646 18672 17651 18728
rect 17585 18667 17651 18672
rect 5498 18528 5818 18529
rect 0 18458 800 18488
rect 5498 18464 5506 18528
rect 5570 18464 5586 18528
rect 5650 18464 5666 18528
rect 5730 18464 5746 18528
rect 5810 18464 5818 18528
rect 5498 18463 5818 18464
rect 14606 18528 14926 18529
rect 14606 18464 14614 18528
rect 14678 18464 14694 18528
rect 14758 18464 14774 18528
rect 14838 18464 14854 18528
rect 14918 18464 14926 18528
rect 14606 18463 14926 18464
rect 23714 18528 24034 18529
rect 23714 18464 23722 18528
rect 23786 18464 23802 18528
rect 23866 18464 23882 18528
rect 23946 18464 23962 18528
rect 24026 18464 24034 18528
rect 23714 18463 24034 18464
rect 1577 18458 1643 18461
rect 0 18456 1643 18458
rect 0 18400 1582 18456
rect 1638 18400 1643 18456
rect 0 18398 1643 18400
rect 0 18368 800 18398
rect 1577 18395 1643 18398
rect 26877 18458 26943 18461
rect 28780 18458 29580 18488
rect 26877 18456 29580 18458
rect 26877 18400 26882 18456
rect 26938 18400 29580 18456
rect 26877 18398 29580 18400
rect 26877 18395 26943 18398
rect 28780 18368 29580 18398
rect 19977 18186 20043 18189
rect 20989 18186 21055 18189
rect 19977 18184 21055 18186
rect 19977 18128 19982 18184
rect 20038 18128 20994 18184
rect 21050 18128 21055 18184
rect 19977 18126 21055 18128
rect 19977 18123 20043 18126
rect 20989 18123 21055 18126
rect 10052 17984 10372 17985
rect 10052 17920 10060 17984
rect 10124 17920 10140 17984
rect 10204 17920 10220 17984
rect 10284 17920 10300 17984
rect 10364 17920 10372 17984
rect 10052 17919 10372 17920
rect 19160 17984 19480 17985
rect 19160 17920 19168 17984
rect 19232 17920 19248 17984
rect 19312 17920 19328 17984
rect 19392 17920 19408 17984
rect 19472 17920 19480 17984
rect 19160 17919 19480 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 25497 17778 25563 17781
rect 28780 17778 29580 17808
rect 25497 17776 29580 17778
rect 25497 17720 25502 17776
rect 25558 17720 29580 17776
rect 25497 17718 29580 17720
rect 25497 17715 25563 17718
rect 28780 17688 29580 17718
rect 14181 17642 14247 17645
rect 16665 17642 16731 17645
rect 14181 17640 16731 17642
rect 14181 17584 14186 17640
rect 14242 17584 16670 17640
rect 16726 17584 16731 17640
rect 14181 17582 16731 17584
rect 14181 17579 14247 17582
rect 16665 17579 16731 17582
rect 5498 17440 5818 17441
rect 5498 17376 5506 17440
rect 5570 17376 5586 17440
rect 5650 17376 5666 17440
rect 5730 17376 5746 17440
rect 5810 17376 5818 17440
rect 5498 17375 5818 17376
rect 14606 17440 14926 17441
rect 14606 17376 14614 17440
rect 14678 17376 14694 17440
rect 14758 17376 14774 17440
rect 14838 17376 14854 17440
rect 14918 17376 14926 17440
rect 14606 17375 14926 17376
rect 23714 17440 24034 17441
rect 23714 17376 23722 17440
rect 23786 17376 23802 17440
rect 23866 17376 23882 17440
rect 23946 17376 23962 17440
rect 24026 17376 24034 17440
rect 23714 17375 24034 17376
rect 9857 17372 9923 17373
rect 9806 17308 9812 17372
rect 9876 17370 9923 17372
rect 9876 17368 9968 17370
rect 9918 17312 9968 17368
rect 9876 17310 9968 17312
rect 9876 17308 9923 17310
rect 9857 17307 9923 17308
rect 19609 17234 19675 17237
rect 21541 17234 21607 17237
rect 19609 17232 21607 17234
rect 19609 17176 19614 17232
rect 19670 17176 21546 17232
rect 21602 17176 21607 17232
rect 19609 17174 21607 17176
rect 19609 17171 19675 17174
rect 21541 17171 21607 17174
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 20713 17098 20779 17101
rect 22737 17098 22803 17101
rect 24945 17098 25011 17101
rect 20713 17096 25011 17098
rect 20713 17040 20718 17096
rect 20774 17040 22742 17096
rect 22798 17040 24950 17096
rect 25006 17040 25011 17096
rect 20713 17038 25011 17040
rect 20713 17035 20779 17038
rect 22737 17035 22803 17038
rect 24945 17035 25011 17038
rect 26141 17098 26207 17101
rect 28780 17098 29580 17128
rect 26141 17096 29580 17098
rect 26141 17040 26146 17096
rect 26202 17040 29580 17096
rect 26141 17038 29580 17040
rect 26141 17035 26207 17038
rect 28780 17008 29580 17038
rect 14089 16962 14155 16965
rect 16021 16962 16087 16965
rect 18045 16962 18111 16965
rect 14089 16960 18111 16962
rect 14089 16904 14094 16960
rect 14150 16904 16026 16960
rect 16082 16904 18050 16960
rect 18106 16904 18111 16960
rect 14089 16902 18111 16904
rect 14089 16899 14155 16902
rect 16021 16899 16087 16902
rect 18045 16899 18111 16902
rect 10052 16896 10372 16897
rect 10052 16832 10060 16896
rect 10124 16832 10140 16896
rect 10204 16832 10220 16896
rect 10284 16832 10300 16896
rect 10364 16832 10372 16896
rect 10052 16831 10372 16832
rect 19160 16896 19480 16897
rect 19160 16832 19168 16896
rect 19232 16832 19248 16896
rect 19312 16832 19328 16896
rect 19392 16832 19408 16896
rect 19472 16832 19480 16896
rect 19160 16831 19480 16832
rect 5498 16352 5818 16353
rect 5498 16288 5506 16352
rect 5570 16288 5586 16352
rect 5650 16288 5666 16352
rect 5730 16288 5746 16352
rect 5810 16288 5818 16352
rect 5498 16287 5818 16288
rect 14606 16352 14926 16353
rect 14606 16288 14614 16352
rect 14678 16288 14694 16352
rect 14758 16288 14774 16352
rect 14838 16288 14854 16352
rect 14918 16288 14926 16352
rect 14606 16287 14926 16288
rect 23714 16352 24034 16353
rect 23714 16288 23722 16352
rect 23786 16288 23802 16352
rect 23866 16288 23882 16352
rect 23946 16288 23962 16352
rect 24026 16288 24034 16352
rect 23714 16287 24034 16288
rect 15193 16282 15259 16285
rect 18229 16282 18295 16285
rect 15193 16280 18295 16282
rect 15193 16224 15198 16280
rect 15254 16224 18234 16280
rect 18290 16224 18295 16280
rect 15193 16222 18295 16224
rect 15193 16219 15259 16222
rect 18229 16219 18295 16222
rect 10910 16084 10916 16148
rect 10980 16146 10986 16148
rect 11053 16146 11119 16149
rect 15929 16146 15995 16149
rect 10980 16144 15995 16146
rect 10980 16088 11058 16144
rect 11114 16088 15934 16144
rect 15990 16088 15995 16144
rect 10980 16086 15995 16088
rect 10980 16084 10986 16086
rect 11053 16083 11119 16086
rect 15929 16083 15995 16086
rect 10052 15808 10372 15809
rect 0 15738 800 15768
rect 10052 15744 10060 15808
rect 10124 15744 10140 15808
rect 10204 15744 10220 15808
rect 10284 15744 10300 15808
rect 10364 15744 10372 15808
rect 10052 15743 10372 15744
rect 19160 15808 19480 15809
rect 19160 15744 19168 15808
rect 19232 15744 19248 15808
rect 19312 15744 19328 15808
rect 19392 15744 19408 15808
rect 19472 15744 19480 15808
rect 19160 15743 19480 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 20805 15738 20871 15741
rect 25129 15738 25195 15741
rect 20805 15736 25195 15738
rect 20805 15680 20810 15736
rect 20866 15680 25134 15736
rect 25190 15680 25195 15736
rect 20805 15678 25195 15680
rect 20805 15675 20871 15678
rect 25129 15675 25195 15678
rect 25589 15738 25655 15741
rect 28780 15738 29580 15768
rect 25589 15736 29580 15738
rect 25589 15680 25594 15736
rect 25650 15680 29580 15736
rect 25589 15678 29580 15680
rect 25589 15675 25655 15678
rect 28780 15648 29580 15678
rect 10869 15466 10935 15469
rect 16297 15466 16363 15469
rect 10869 15464 16363 15466
rect 10869 15408 10874 15464
rect 10930 15408 16302 15464
rect 16358 15408 16363 15464
rect 10869 15406 16363 15408
rect 10869 15403 10935 15406
rect 16297 15403 16363 15406
rect 19885 15330 19951 15333
rect 22093 15330 22159 15333
rect 19885 15328 22159 15330
rect 19885 15272 19890 15328
rect 19946 15272 22098 15328
rect 22154 15272 22159 15328
rect 19885 15270 22159 15272
rect 19885 15267 19951 15270
rect 22093 15267 22159 15270
rect 5498 15264 5818 15265
rect 5498 15200 5506 15264
rect 5570 15200 5586 15264
rect 5650 15200 5666 15264
rect 5730 15200 5746 15264
rect 5810 15200 5818 15264
rect 5498 15199 5818 15200
rect 14606 15264 14926 15265
rect 14606 15200 14614 15264
rect 14678 15200 14694 15264
rect 14758 15200 14774 15264
rect 14838 15200 14854 15264
rect 14918 15200 14926 15264
rect 14606 15199 14926 15200
rect 23714 15264 24034 15265
rect 23714 15200 23722 15264
rect 23786 15200 23802 15264
rect 23866 15200 23882 15264
rect 23946 15200 23962 15264
rect 24026 15200 24034 15264
rect 23714 15199 24034 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 13077 15058 13143 15061
rect 18965 15058 19031 15061
rect 13077 15056 19031 15058
rect 13077 15000 13082 15056
rect 13138 15000 18970 15056
rect 19026 15000 19031 15056
rect 13077 14998 19031 15000
rect 13077 14995 13143 14998
rect 18965 14995 19031 14998
rect 26877 15058 26943 15061
rect 28780 15058 29580 15088
rect 26877 15056 29580 15058
rect 26877 15000 26882 15056
rect 26938 15000 29580 15056
rect 26877 14998 29580 15000
rect 26877 14995 26943 14998
rect 28780 14968 29580 14998
rect 9121 14922 9187 14925
rect 9581 14922 9647 14925
rect 14089 14922 14155 14925
rect 9121 14920 14155 14922
rect 9121 14864 9126 14920
rect 9182 14864 9586 14920
rect 9642 14864 14094 14920
rect 14150 14864 14155 14920
rect 9121 14862 14155 14864
rect 9121 14859 9187 14862
rect 9581 14859 9647 14862
rect 14089 14859 14155 14862
rect 14825 14922 14891 14925
rect 15561 14922 15627 14925
rect 19701 14922 19767 14925
rect 14825 14920 19767 14922
rect 14825 14864 14830 14920
rect 14886 14864 15566 14920
rect 15622 14864 19706 14920
rect 19762 14864 19767 14920
rect 14825 14862 19767 14864
rect 14825 14859 14891 14862
rect 15561 14859 15627 14862
rect 19701 14859 19767 14862
rect 21357 14922 21423 14925
rect 22185 14922 22251 14925
rect 24209 14922 24275 14925
rect 21357 14920 24275 14922
rect 21357 14864 21362 14920
rect 21418 14864 22190 14920
rect 22246 14864 24214 14920
rect 24270 14864 24275 14920
rect 21357 14862 24275 14864
rect 21357 14859 21423 14862
rect 22185 14859 22251 14862
rect 24209 14859 24275 14862
rect 14917 14786 14983 14789
rect 15193 14786 15259 14789
rect 18505 14786 18571 14789
rect 14917 14784 15259 14786
rect 14917 14728 14922 14784
rect 14978 14728 15198 14784
rect 15254 14728 15259 14784
rect 14917 14726 15259 14728
rect 14917 14723 14983 14726
rect 15193 14723 15259 14726
rect 15334 14784 18571 14786
rect 15334 14728 18510 14784
rect 18566 14728 18571 14784
rect 15334 14726 18571 14728
rect 10052 14720 10372 14721
rect 10052 14656 10060 14720
rect 10124 14656 10140 14720
rect 10204 14656 10220 14720
rect 10284 14656 10300 14720
rect 10364 14656 10372 14720
rect 10052 14655 10372 14656
rect 10777 14650 10843 14653
rect 15334 14650 15394 14726
rect 18505 14723 18571 14726
rect 19160 14720 19480 14721
rect 19160 14656 19168 14720
rect 19232 14656 19248 14720
rect 19312 14656 19328 14720
rect 19392 14656 19408 14720
rect 19472 14656 19480 14720
rect 19160 14655 19480 14656
rect 10777 14648 15394 14650
rect 10777 14592 10782 14648
rect 10838 14592 15394 14648
rect 10777 14590 15394 14592
rect 17585 14650 17651 14653
rect 17953 14650 18019 14653
rect 17585 14648 18019 14650
rect 17585 14592 17590 14648
rect 17646 14592 17958 14648
rect 18014 14592 18019 14648
rect 17585 14590 18019 14592
rect 10777 14587 10843 14590
rect 17585 14587 17651 14590
rect 17953 14587 18019 14590
rect 1853 14514 1919 14517
rect 9121 14514 9187 14517
rect 1853 14512 9187 14514
rect 1853 14456 1858 14512
rect 1914 14456 9126 14512
rect 9182 14456 9187 14512
rect 1853 14454 9187 14456
rect 1853 14451 1919 14454
rect 9121 14451 9187 14454
rect 14181 14514 14247 14517
rect 17217 14514 17283 14517
rect 18505 14514 18571 14517
rect 14181 14512 18571 14514
rect 14181 14456 14186 14512
rect 14242 14456 17222 14512
rect 17278 14456 18510 14512
rect 18566 14456 18571 14512
rect 14181 14454 18571 14456
rect 14181 14451 14247 14454
rect 17217 14451 17283 14454
rect 18505 14451 18571 14454
rect 0 14378 800 14408
rect 2037 14378 2103 14381
rect 0 14376 2103 14378
rect 0 14320 2042 14376
rect 2098 14320 2103 14376
rect 0 14318 2103 14320
rect 0 14288 800 14318
rect 2037 14315 2103 14318
rect 7833 14378 7899 14381
rect 8569 14378 8635 14381
rect 7833 14376 8635 14378
rect 7833 14320 7838 14376
rect 7894 14320 8574 14376
rect 8630 14320 8635 14376
rect 7833 14318 8635 14320
rect 7833 14315 7899 14318
rect 8569 14315 8635 14318
rect 10317 14378 10383 14381
rect 14733 14378 14799 14381
rect 10317 14376 14799 14378
rect 10317 14320 10322 14376
rect 10378 14320 14738 14376
rect 14794 14320 14799 14376
rect 10317 14318 14799 14320
rect 10317 14315 10383 14318
rect 14733 14315 14799 14318
rect 26141 14378 26207 14381
rect 28780 14378 29580 14408
rect 26141 14376 29580 14378
rect 26141 14320 26146 14376
rect 26202 14320 29580 14376
rect 26141 14318 29580 14320
rect 26141 14315 26207 14318
rect 28780 14288 29580 14318
rect 5498 14176 5818 14177
rect 5498 14112 5506 14176
rect 5570 14112 5586 14176
rect 5650 14112 5666 14176
rect 5730 14112 5746 14176
rect 5810 14112 5818 14176
rect 5498 14111 5818 14112
rect 14606 14176 14926 14177
rect 14606 14112 14614 14176
rect 14678 14112 14694 14176
rect 14758 14112 14774 14176
rect 14838 14112 14854 14176
rect 14918 14112 14926 14176
rect 14606 14111 14926 14112
rect 23714 14176 24034 14177
rect 23714 14112 23722 14176
rect 23786 14112 23802 14176
rect 23866 14112 23882 14176
rect 23946 14112 23962 14176
rect 24026 14112 24034 14176
rect 23714 14111 24034 14112
rect 10777 13970 10843 13973
rect 12157 13970 12223 13973
rect 10777 13968 12223 13970
rect 10777 13912 10782 13968
rect 10838 13912 12162 13968
rect 12218 13912 12223 13968
rect 10777 13910 12223 13912
rect 10777 13907 10843 13910
rect 12157 13907 12223 13910
rect 17953 13970 18019 13973
rect 18229 13970 18295 13973
rect 17953 13968 18295 13970
rect 17953 13912 17958 13968
rect 18014 13912 18234 13968
rect 18290 13912 18295 13968
rect 17953 13910 18295 13912
rect 17953 13907 18019 13910
rect 18229 13907 18295 13910
rect 9765 13834 9831 13837
rect 10593 13834 10659 13837
rect 16205 13834 16271 13837
rect 9765 13832 16271 13834
rect 9765 13776 9770 13832
rect 9826 13776 10598 13832
rect 10654 13776 16210 13832
rect 16266 13776 16271 13832
rect 9765 13774 16271 13776
rect 9765 13771 9831 13774
rect 10593 13771 10659 13774
rect 16205 13771 16271 13774
rect 10052 13632 10372 13633
rect 10052 13568 10060 13632
rect 10124 13568 10140 13632
rect 10204 13568 10220 13632
rect 10284 13568 10300 13632
rect 10364 13568 10372 13632
rect 10052 13567 10372 13568
rect 19160 13632 19480 13633
rect 19160 13568 19168 13632
rect 19232 13568 19248 13632
rect 19312 13568 19328 13632
rect 19392 13568 19408 13632
rect 19472 13568 19480 13632
rect 19160 13567 19480 13568
rect 5498 13088 5818 13089
rect 0 13018 800 13048
rect 5498 13024 5506 13088
rect 5570 13024 5586 13088
rect 5650 13024 5666 13088
rect 5730 13024 5746 13088
rect 5810 13024 5818 13088
rect 5498 13023 5818 13024
rect 14606 13088 14926 13089
rect 14606 13024 14614 13088
rect 14678 13024 14694 13088
rect 14758 13024 14774 13088
rect 14838 13024 14854 13088
rect 14918 13024 14926 13088
rect 14606 13023 14926 13024
rect 23714 13088 24034 13089
rect 23714 13024 23722 13088
rect 23786 13024 23802 13088
rect 23866 13024 23882 13088
rect 23946 13024 23962 13088
rect 24026 13024 24034 13088
rect 23714 13023 24034 13024
rect 1393 13018 1459 13021
rect 0 13016 1459 13018
rect 0 12960 1398 13016
rect 1454 12960 1459 13016
rect 0 12958 1459 12960
rect 0 12928 800 12958
rect 1393 12955 1459 12958
rect 27797 13018 27863 13021
rect 28780 13018 29580 13048
rect 27797 13016 29580 13018
rect 27797 12960 27802 13016
rect 27858 12960 29580 13016
rect 27797 12958 29580 12960
rect 27797 12955 27863 12958
rect 28780 12928 29580 12958
rect 7097 12882 7163 12885
rect 7925 12882 7991 12885
rect 7097 12880 7991 12882
rect 7097 12824 7102 12880
rect 7158 12824 7930 12880
rect 7986 12824 7991 12880
rect 7097 12822 7991 12824
rect 7097 12819 7163 12822
rect 7925 12819 7991 12822
rect 15745 12882 15811 12885
rect 18229 12882 18295 12885
rect 15745 12880 18295 12882
rect 15745 12824 15750 12880
rect 15806 12824 18234 12880
rect 18290 12824 18295 12880
rect 15745 12822 18295 12824
rect 15745 12819 15811 12822
rect 18229 12819 18295 12822
rect 4889 12746 4955 12749
rect 9581 12746 9647 12749
rect 4889 12744 9647 12746
rect 4889 12688 4894 12744
rect 4950 12688 9586 12744
rect 9642 12688 9647 12744
rect 4889 12686 9647 12688
rect 4889 12683 4955 12686
rect 9581 12683 9647 12686
rect 15929 12610 15995 12613
rect 18321 12610 18387 12613
rect 15929 12608 18387 12610
rect 15929 12552 15934 12608
rect 15990 12552 18326 12608
rect 18382 12552 18387 12608
rect 15929 12550 18387 12552
rect 15929 12547 15995 12550
rect 18321 12547 18387 12550
rect 10052 12544 10372 12545
rect 10052 12480 10060 12544
rect 10124 12480 10140 12544
rect 10204 12480 10220 12544
rect 10284 12480 10300 12544
rect 10364 12480 10372 12544
rect 10052 12479 10372 12480
rect 19160 12544 19480 12545
rect 19160 12480 19168 12544
rect 19232 12480 19248 12544
rect 19312 12480 19328 12544
rect 19392 12480 19408 12544
rect 19472 12480 19480 12544
rect 19160 12479 19480 12480
rect 15837 12474 15903 12477
rect 18965 12474 19031 12477
rect 15837 12472 19031 12474
rect 15837 12416 15842 12472
rect 15898 12416 18970 12472
rect 19026 12416 19031 12472
rect 15837 12414 19031 12416
rect 15837 12411 15903 12414
rect 18965 12411 19031 12414
rect 0 12338 800 12368
rect 2037 12338 2103 12341
rect 0 12336 2103 12338
rect 0 12280 2042 12336
rect 2098 12280 2103 12336
rect 0 12278 2103 12280
rect 0 12248 800 12278
rect 2037 12275 2103 12278
rect 27705 12338 27771 12341
rect 28780 12338 29580 12368
rect 27705 12336 29580 12338
rect 27705 12280 27710 12336
rect 27766 12280 29580 12336
rect 27705 12278 29580 12280
rect 27705 12275 27771 12278
rect 28780 12248 29580 12278
rect 7281 12202 7347 12205
rect 7833 12202 7899 12205
rect 7281 12200 7899 12202
rect 7281 12144 7286 12200
rect 7342 12144 7838 12200
rect 7894 12144 7899 12200
rect 7281 12142 7899 12144
rect 7281 12139 7347 12142
rect 7833 12139 7899 12142
rect 5498 12000 5818 12001
rect 5498 11936 5506 12000
rect 5570 11936 5586 12000
rect 5650 11936 5666 12000
rect 5730 11936 5746 12000
rect 5810 11936 5818 12000
rect 5498 11935 5818 11936
rect 14606 12000 14926 12001
rect 14606 11936 14614 12000
rect 14678 11936 14694 12000
rect 14758 11936 14774 12000
rect 14838 11936 14854 12000
rect 14918 11936 14926 12000
rect 14606 11935 14926 11936
rect 23714 12000 24034 12001
rect 23714 11936 23722 12000
rect 23786 11936 23802 12000
rect 23866 11936 23882 12000
rect 23946 11936 23962 12000
rect 24026 11936 24034 12000
rect 23714 11935 24034 11936
rect 16849 11930 16915 11933
rect 17309 11930 17375 11933
rect 16849 11928 17375 11930
rect 16849 11872 16854 11928
rect 16910 11872 17314 11928
rect 17370 11872 17375 11928
rect 16849 11870 17375 11872
rect 16849 11867 16915 11870
rect 17309 11867 17375 11870
rect 20805 11794 20871 11797
rect 21173 11794 21239 11797
rect 22001 11794 22067 11797
rect 24209 11794 24275 11797
rect 20805 11792 24275 11794
rect 20805 11736 20810 11792
rect 20866 11736 21178 11792
rect 21234 11736 22006 11792
rect 22062 11736 24214 11792
rect 24270 11736 24275 11792
rect 20805 11734 24275 11736
rect 20805 11731 20871 11734
rect 21173 11731 21239 11734
rect 22001 11731 22067 11734
rect 24209 11731 24275 11734
rect 0 11658 800 11688
rect 1669 11658 1735 11661
rect 0 11656 1735 11658
rect 0 11600 1674 11656
rect 1730 11600 1735 11656
rect 0 11598 1735 11600
rect 0 11568 800 11598
rect 1669 11595 1735 11598
rect 26877 11658 26943 11661
rect 28780 11658 29580 11688
rect 26877 11656 29580 11658
rect 26877 11600 26882 11656
rect 26938 11600 29580 11656
rect 26877 11598 29580 11600
rect 26877 11595 26943 11598
rect 28780 11568 29580 11598
rect 10052 11456 10372 11457
rect 10052 11392 10060 11456
rect 10124 11392 10140 11456
rect 10204 11392 10220 11456
rect 10284 11392 10300 11456
rect 10364 11392 10372 11456
rect 10052 11391 10372 11392
rect 19160 11456 19480 11457
rect 19160 11392 19168 11456
rect 19232 11392 19248 11456
rect 19312 11392 19328 11456
rect 19392 11392 19408 11456
rect 19472 11392 19480 11456
rect 19160 11391 19480 11392
rect 21265 11250 21331 11253
rect 23197 11250 23263 11253
rect 23749 11250 23815 11253
rect 21265 11248 23815 11250
rect 21265 11192 21270 11248
rect 21326 11192 23202 11248
rect 23258 11192 23754 11248
rect 23810 11192 23815 11248
rect 21265 11190 23815 11192
rect 21265 11187 21331 11190
rect 23197 11187 23263 11190
rect 23749 11187 23815 11190
rect 9029 11114 9095 11117
rect 10685 11114 10751 11117
rect 10910 11114 10916 11116
rect 9029 11112 10916 11114
rect 9029 11056 9034 11112
rect 9090 11056 10690 11112
rect 10746 11056 10916 11112
rect 9029 11054 10916 11056
rect 9029 11051 9095 11054
rect 10685 11051 10751 11054
rect 10910 11052 10916 11054
rect 10980 11052 10986 11116
rect 8477 10978 8543 10981
rect 10409 10978 10475 10981
rect 12157 10978 12223 10981
rect 8477 10976 12223 10978
rect 8477 10920 8482 10976
rect 8538 10920 10414 10976
rect 10470 10920 12162 10976
rect 12218 10920 12223 10976
rect 8477 10918 12223 10920
rect 8477 10915 8543 10918
rect 10409 10915 10475 10918
rect 12157 10915 12223 10918
rect 5498 10912 5818 10913
rect 5498 10848 5506 10912
rect 5570 10848 5586 10912
rect 5650 10848 5666 10912
rect 5730 10848 5746 10912
rect 5810 10848 5818 10912
rect 5498 10847 5818 10848
rect 14606 10912 14926 10913
rect 14606 10848 14614 10912
rect 14678 10848 14694 10912
rect 14758 10848 14774 10912
rect 14838 10848 14854 10912
rect 14918 10848 14926 10912
rect 14606 10847 14926 10848
rect 23714 10912 24034 10913
rect 23714 10848 23722 10912
rect 23786 10848 23802 10912
rect 23866 10848 23882 10912
rect 23946 10848 23962 10912
rect 24026 10848 24034 10912
rect 23714 10847 24034 10848
rect 10052 10368 10372 10369
rect 0 10298 800 10328
rect 10052 10304 10060 10368
rect 10124 10304 10140 10368
rect 10204 10304 10220 10368
rect 10284 10304 10300 10368
rect 10364 10304 10372 10368
rect 10052 10303 10372 10304
rect 19160 10368 19480 10369
rect 19160 10304 19168 10368
rect 19232 10304 19248 10368
rect 19312 10304 19328 10368
rect 19392 10304 19408 10368
rect 19472 10304 19480 10368
rect 19160 10303 19480 10304
rect 1945 10298 2011 10301
rect 0 10296 2011 10298
rect 0 10240 1950 10296
rect 2006 10240 2011 10296
rect 0 10238 2011 10240
rect 0 10208 800 10238
rect 1945 10235 2011 10238
rect 26785 10298 26851 10301
rect 28780 10298 29580 10328
rect 26785 10296 29580 10298
rect 26785 10240 26790 10296
rect 26846 10240 29580 10296
rect 26785 10238 29580 10240
rect 26785 10235 26851 10238
rect 28780 10208 29580 10238
rect 5498 9824 5818 9825
rect 5498 9760 5506 9824
rect 5570 9760 5586 9824
rect 5650 9760 5666 9824
rect 5730 9760 5746 9824
rect 5810 9760 5818 9824
rect 5498 9759 5818 9760
rect 14606 9824 14926 9825
rect 14606 9760 14614 9824
rect 14678 9760 14694 9824
rect 14758 9760 14774 9824
rect 14838 9760 14854 9824
rect 14918 9760 14926 9824
rect 14606 9759 14926 9760
rect 23714 9824 24034 9825
rect 23714 9760 23722 9824
rect 23786 9760 23802 9824
rect 23866 9760 23882 9824
rect 23946 9760 23962 9824
rect 24026 9760 24034 9824
rect 23714 9759 24034 9760
rect 12157 9754 12223 9757
rect 13905 9754 13971 9757
rect 12157 9752 13971 9754
rect 12157 9696 12162 9752
rect 12218 9696 13910 9752
rect 13966 9696 13971 9752
rect 12157 9694 13971 9696
rect 12157 9691 12223 9694
rect 13905 9691 13971 9694
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 20897 9618 20963 9621
rect 22001 9618 22067 9621
rect 20897 9616 22067 9618
rect 20897 9560 20902 9616
rect 20958 9560 22006 9616
rect 22062 9560 22067 9616
rect 20897 9558 22067 9560
rect 20897 9555 20963 9558
rect 22001 9555 22067 9558
rect 26693 9618 26759 9621
rect 28780 9618 29580 9648
rect 26693 9616 29580 9618
rect 26693 9560 26698 9616
rect 26754 9560 29580 9616
rect 26693 9558 29580 9560
rect 26693 9555 26759 9558
rect 28780 9528 29580 9558
rect 9806 9420 9812 9484
rect 9876 9482 9882 9484
rect 10317 9482 10383 9485
rect 9876 9480 10383 9482
rect 9876 9424 10322 9480
rect 10378 9424 10383 9480
rect 9876 9422 10383 9424
rect 9876 9420 9882 9422
rect 10317 9419 10383 9422
rect 10052 9280 10372 9281
rect 10052 9216 10060 9280
rect 10124 9216 10140 9280
rect 10204 9216 10220 9280
rect 10284 9216 10300 9280
rect 10364 9216 10372 9280
rect 10052 9215 10372 9216
rect 19160 9280 19480 9281
rect 19160 9216 19168 9280
rect 19232 9216 19248 9280
rect 19312 9216 19328 9280
rect 19392 9216 19408 9280
rect 19472 9216 19480 9280
rect 19160 9215 19480 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 19885 8938 19951 8941
rect 27521 8938 27587 8941
rect 19885 8936 27587 8938
rect 19885 8880 19890 8936
rect 19946 8880 27526 8936
rect 27582 8880 27587 8936
rect 19885 8878 27587 8880
rect 19885 8875 19951 8878
rect 27521 8875 27587 8878
rect 27705 8938 27771 8941
rect 28780 8938 29580 8968
rect 27705 8936 29580 8938
rect 27705 8880 27710 8936
rect 27766 8880 29580 8936
rect 27705 8878 29580 8880
rect 27705 8875 27771 8878
rect 28780 8848 29580 8878
rect 5498 8736 5818 8737
rect 5498 8672 5506 8736
rect 5570 8672 5586 8736
rect 5650 8672 5666 8736
rect 5730 8672 5746 8736
rect 5810 8672 5818 8736
rect 5498 8671 5818 8672
rect 14606 8736 14926 8737
rect 14606 8672 14614 8736
rect 14678 8672 14694 8736
rect 14758 8672 14774 8736
rect 14838 8672 14854 8736
rect 14918 8672 14926 8736
rect 14606 8671 14926 8672
rect 23714 8736 24034 8737
rect 23714 8672 23722 8736
rect 23786 8672 23802 8736
rect 23866 8672 23882 8736
rect 23946 8672 23962 8736
rect 24026 8672 24034 8736
rect 23714 8671 24034 8672
rect 14181 8530 14247 8533
rect 18965 8530 19031 8533
rect 14181 8528 19031 8530
rect 14181 8472 14186 8528
rect 14242 8472 18970 8528
rect 19026 8472 19031 8528
rect 14181 8470 19031 8472
rect 14181 8467 14247 8470
rect 18965 8467 19031 8470
rect 9765 8394 9831 8397
rect 13537 8394 13603 8397
rect 9765 8392 13603 8394
rect 9765 8336 9770 8392
rect 9826 8336 13542 8392
rect 13598 8336 13603 8392
rect 9765 8334 13603 8336
rect 9765 8331 9831 8334
rect 13537 8331 13603 8334
rect 10052 8192 10372 8193
rect 10052 8128 10060 8192
rect 10124 8128 10140 8192
rect 10204 8128 10220 8192
rect 10284 8128 10300 8192
rect 10364 8128 10372 8192
rect 10052 8127 10372 8128
rect 19160 8192 19480 8193
rect 19160 8128 19168 8192
rect 19232 8128 19248 8192
rect 19312 8128 19328 8192
rect 19392 8128 19408 8192
rect 19472 8128 19480 8192
rect 19160 8127 19480 8128
rect 4429 7986 4495 7989
rect 6085 7986 6151 7989
rect 4429 7984 6151 7986
rect 4429 7928 4434 7984
rect 4490 7928 6090 7984
rect 6146 7928 6151 7984
rect 4429 7926 6151 7928
rect 4429 7923 4495 7926
rect 6085 7923 6151 7926
rect 20897 7986 20963 7989
rect 23013 7986 23079 7989
rect 20897 7984 23079 7986
rect 20897 7928 20902 7984
rect 20958 7928 23018 7984
rect 23074 7928 23079 7984
rect 20897 7926 23079 7928
rect 20897 7923 20963 7926
rect 23013 7923 23079 7926
rect 20253 7850 20319 7853
rect 22829 7850 22895 7853
rect 20253 7848 22895 7850
rect 20253 7792 20258 7848
rect 20314 7792 22834 7848
rect 22890 7792 22895 7848
rect 20253 7790 22895 7792
rect 20253 7787 20319 7790
rect 22829 7787 22895 7790
rect 5498 7648 5818 7649
rect 0 7578 800 7608
rect 5498 7584 5506 7648
rect 5570 7584 5586 7648
rect 5650 7584 5666 7648
rect 5730 7584 5746 7648
rect 5810 7584 5818 7648
rect 5498 7583 5818 7584
rect 14606 7648 14926 7649
rect 14606 7584 14614 7648
rect 14678 7584 14694 7648
rect 14758 7584 14774 7648
rect 14838 7584 14854 7648
rect 14918 7584 14926 7648
rect 14606 7583 14926 7584
rect 23714 7648 24034 7649
rect 23714 7584 23722 7648
rect 23786 7584 23802 7648
rect 23866 7584 23882 7648
rect 23946 7584 23962 7648
rect 24026 7584 24034 7648
rect 23714 7583 24034 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 26693 7578 26759 7581
rect 28780 7578 29580 7608
rect 26693 7576 29580 7578
rect 26693 7520 26698 7576
rect 26754 7520 29580 7576
rect 26693 7518 29580 7520
rect 26693 7515 26759 7518
rect 28780 7488 29580 7518
rect 10052 7104 10372 7105
rect 10052 7040 10060 7104
rect 10124 7040 10140 7104
rect 10204 7040 10220 7104
rect 10284 7040 10300 7104
rect 10364 7040 10372 7104
rect 10052 7039 10372 7040
rect 19160 7104 19480 7105
rect 19160 7040 19168 7104
rect 19232 7040 19248 7104
rect 19312 7040 19328 7104
rect 19392 7040 19408 7104
rect 19472 7040 19480 7104
rect 19160 7039 19480 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 26141 6898 26207 6901
rect 28780 6898 29580 6928
rect 26141 6896 29580 6898
rect 26141 6840 26146 6896
rect 26202 6840 29580 6896
rect 26141 6838 29580 6840
rect 26141 6835 26207 6838
rect 28780 6808 29580 6838
rect 5498 6560 5818 6561
rect 5498 6496 5506 6560
rect 5570 6496 5586 6560
rect 5650 6496 5666 6560
rect 5730 6496 5746 6560
rect 5810 6496 5818 6560
rect 5498 6495 5818 6496
rect 14606 6560 14926 6561
rect 14606 6496 14614 6560
rect 14678 6496 14694 6560
rect 14758 6496 14774 6560
rect 14838 6496 14854 6560
rect 14918 6496 14926 6560
rect 14606 6495 14926 6496
rect 23714 6560 24034 6561
rect 23714 6496 23722 6560
rect 23786 6496 23802 6560
rect 23866 6496 23882 6560
rect 23946 6496 23962 6560
rect 24026 6496 24034 6560
rect 23714 6495 24034 6496
rect 6269 6354 6335 6357
rect 8477 6354 8543 6357
rect 6269 6352 8543 6354
rect 6269 6296 6274 6352
rect 6330 6296 8482 6352
rect 8538 6296 8543 6352
rect 6269 6294 8543 6296
rect 6269 6291 6335 6294
rect 8477 6291 8543 6294
rect 10133 6354 10199 6357
rect 17677 6354 17743 6357
rect 10133 6352 17743 6354
rect 10133 6296 10138 6352
rect 10194 6296 17682 6352
rect 17738 6296 17743 6352
rect 10133 6294 17743 6296
rect 10133 6291 10199 6294
rect 17677 6291 17743 6294
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 12249 6218 12315 6221
rect 13997 6218 14063 6221
rect 12249 6216 14063 6218
rect 12249 6160 12254 6216
rect 12310 6160 14002 6216
rect 14058 6160 14063 6216
rect 12249 6158 14063 6160
rect 12249 6155 12315 6158
rect 13997 6155 14063 6158
rect 23105 6218 23171 6221
rect 24761 6218 24827 6221
rect 23105 6216 24827 6218
rect 23105 6160 23110 6216
rect 23166 6160 24766 6216
rect 24822 6160 24827 6216
rect 23105 6158 24827 6160
rect 23105 6155 23171 6158
rect 24761 6155 24827 6158
rect 27705 6218 27771 6221
rect 28780 6218 29580 6248
rect 27705 6216 29580 6218
rect 27705 6160 27710 6216
rect 27766 6160 29580 6216
rect 27705 6158 29580 6160
rect 27705 6155 27771 6158
rect 28780 6128 29580 6158
rect 10052 6016 10372 6017
rect 10052 5952 10060 6016
rect 10124 5952 10140 6016
rect 10204 5952 10220 6016
rect 10284 5952 10300 6016
rect 10364 5952 10372 6016
rect 10052 5951 10372 5952
rect 19160 6016 19480 6017
rect 19160 5952 19168 6016
rect 19232 5952 19248 6016
rect 19312 5952 19328 6016
rect 19392 5952 19408 6016
rect 19472 5952 19480 6016
rect 19160 5951 19480 5952
rect 8569 5810 8635 5813
rect 9857 5810 9923 5813
rect 8569 5808 9923 5810
rect 8569 5752 8574 5808
rect 8630 5752 9862 5808
rect 9918 5752 9923 5808
rect 8569 5750 9923 5752
rect 8569 5747 8635 5750
rect 9857 5747 9923 5750
rect 5498 5472 5818 5473
rect 5498 5408 5506 5472
rect 5570 5408 5586 5472
rect 5650 5408 5666 5472
rect 5730 5408 5746 5472
rect 5810 5408 5818 5472
rect 5498 5407 5818 5408
rect 14606 5472 14926 5473
rect 14606 5408 14614 5472
rect 14678 5408 14694 5472
rect 14758 5408 14774 5472
rect 14838 5408 14854 5472
rect 14918 5408 14926 5472
rect 14606 5407 14926 5408
rect 23714 5472 24034 5473
rect 23714 5408 23722 5472
rect 23786 5408 23802 5472
rect 23866 5408 23882 5472
rect 23946 5408 23962 5472
rect 24026 5408 24034 5472
rect 23714 5407 24034 5408
rect 10052 4928 10372 4929
rect 0 4858 800 4888
rect 10052 4864 10060 4928
rect 10124 4864 10140 4928
rect 10204 4864 10220 4928
rect 10284 4864 10300 4928
rect 10364 4864 10372 4928
rect 10052 4863 10372 4864
rect 19160 4928 19480 4929
rect 19160 4864 19168 4928
rect 19232 4864 19248 4928
rect 19312 4864 19328 4928
rect 19392 4864 19408 4928
rect 19472 4864 19480 4928
rect 19160 4863 19480 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 27521 4858 27587 4861
rect 28780 4858 29580 4888
rect 27521 4856 29580 4858
rect 27521 4800 27526 4856
rect 27582 4800 29580 4856
rect 27521 4798 29580 4800
rect 27521 4795 27587 4798
rect 28780 4768 29580 4798
rect 10685 4722 10751 4725
rect 11697 4722 11763 4725
rect 13261 4722 13327 4725
rect 10685 4720 13327 4722
rect 10685 4664 10690 4720
rect 10746 4664 11702 4720
rect 11758 4664 13266 4720
rect 13322 4664 13327 4720
rect 10685 4662 13327 4664
rect 10685 4659 10751 4662
rect 11697 4659 11763 4662
rect 13261 4659 13327 4662
rect 19701 4722 19767 4725
rect 20621 4722 20687 4725
rect 19701 4720 20687 4722
rect 19701 4664 19706 4720
rect 19762 4664 20626 4720
rect 20682 4664 20687 4720
rect 19701 4662 20687 4664
rect 19701 4659 19767 4662
rect 20621 4659 20687 4662
rect 17217 4450 17283 4453
rect 23013 4450 23079 4453
rect 17217 4448 23079 4450
rect 17217 4392 17222 4448
rect 17278 4392 23018 4448
rect 23074 4392 23079 4448
rect 17217 4390 23079 4392
rect 17217 4387 17283 4390
rect 23013 4387 23079 4390
rect 5498 4384 5818 4385
rect 5498 4320 5506 4384
rect 5570 4320 5586 4384
rect 5650 4320 5666 4384
rect 5730 4320 5746 4384
rect 5810 4320 5818 4384
rect 5498 4319 5818 4320
rect 14606 4384 14926 4385
rect 14606 4320 14614 4384
rect 14678 4320 14694 4384
rect 14758 4320 14774 4384
rect 14838 4320 14854 4384
rect 14918 4320 14926 4384
rect 14606 4319 14926 4320
rect 23714 4384 24034 4385
rect 23714 4320 23722 4384
rect 23786 4320 23802 4384
rect 23866 4320 23882 4384
rect 23946 4320 23962 4384
rect 24026 4320 24034 4384
rect 23714 4319 24034 4320
rect 0 4178 800 4208
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4088 800 4118
rect 2773 4115 2839 4118
rect 12525 4178 12591 4181
rect 20713 4178 20779 4181
rect 12525 4176 20779 4178
rect 12525 4120 12530 4176
rect 12586 4120 20718 4176
rect 20774 4120 20779 4176
rect 12525 4118 20779 4120
rect 12525 4115 12591 4118
rect 20713 4115 20779 4118
rect 26785 4178 26851 4181
rect 28780 4178 29580 4208
rect 26785 4176 29580 4178
rect 26785 4120 26790 4176
rect 26846 4120 29580 4176
rect 26785 4118 29580 4120
rect 26785 4115 26851 4118
rect 28780 4088 29580 4118
rect 12341 4042 12407 4045
rect 13169 4042 13235 4045
rect 12341 4040 13235 4042
rect 12341 3984 12346 4040
rect 12402 3984 13174 4040
rect 13230 3984 13235 4040
rect 12341 3982 13235 3984
rect 12341 3979 12407 3982
rect 13169 3979 13235 3982
rect 16113 4042 16179 4045
rect 23933 4042 23999 4045
rect 16113 4040 23999 4042
rect 16113 3984 16118 4040
rect 16174 3984 23938 4040
rect 23994 3984 23999 4040
rect 16113 3982 23999 3984
rect 16113 3979 16179 3982
rect 23933 3979 23999 3982
rect 26141 4042 26207 4045
rect 26366 4042 26372 4044
rect 26141 4040 26372 4042
rect 26141 3984 26146 4040
rect 26202 3984 26372 4040
rect 26141 3982 26372 3984
rect 26141 3979 26207 3982
rect 26366 3980 26372 3982
rect 26436 3980 26442 4044
rect 10052 3840 10372 3841
rect 10052 3776 10060 3840
rect 10124 3776 10140 3840
rect 10204 3776 10220 3840
rect 10284 3776 10300 3840
rect 10364 3776 10372 3840
rect 10052 3775 10372 3776
rect 19160 3840 19480 3841
rect 19160 3776 19168 3840
rect 19232 3776 19248 3840
rect 19312 3776 19328 3840
rect 19392 3776 19408 3840
rect 19472 3776 19480 3840
rect 19160 3775 19480 3776
rect 12985 3770 13051 3773
rect 20253 3770 20319 3773
rect 24393 3770 24459 3773
rect 12985 3768 13186 3770
rect 12985 3712 12990 3768
rect 13046 3712 13186 3768
rect 12985 3710 13186 3712
rect 12985 3707 13051 3710
rect 9673 3634 9739 3637
rect 12893 3634 12959 3637
rect 9673 3632 12959 3634
rect 9673 3576 9678 3632
rect 9734 3576 12898 3632
rect 12954 3576 12959 3632
rect 9673 3574 12959 3576
rect 13126 3634 13186 3710
rect 20253 3768 24459 3770
rect 20253 3712 20258 3768
rect 20314 3712 24398 3768
rect 24454 3712 24459 3768
rect 20253 3710 24459 3712
rect 20253 3707 20319 3710
rect 24393 3707 24459 3710
rect 19149 3634 19215 3637
rect 13126 3632 19215 3634
rect 13126 3576 19154 3632
rect 19210 3576 19215 3632
rect 13126 3574 19215 3576
rect 9673 3571 9739 3574
rect 12893 3571 12959 3574
rect 19149 3571 19215 3574
rect 0 3498 800 3528
rect 3141 3498 3207 3501
rect 0 3496 3207 3498
rect 0 3440 3146 3496
rect 3202 3440 3207 3496
rect 0 3438 3207 3440
rect 0 3408 800 3438
rect 3141 3435 3207 3438
rect 15469 3498 15535 3501
rect 18505 3498 18571 3501
rect 15469 3496 18571 3498
rect 15469 3440 15474 3496
rect 15530 3440 18510 3496
rect 18566 3440 18571 3496
rect 15469 3438 18571 3440
rect 15469 3435 15535 3438
rect 18505 3435 18571 3438
rect 26877 3498 26943 3501
rect 28780 3498 29580 3528
rect 26877 3496 29580 3498
rect 26877 3440 26882 3496
rect 26938 3440 29580 3496
rect 26877 3438 29580 3440
rect 26877 3435 26943 3438
rect 28780 3408 29580 3438
rect 5498 3296 5818 3297
rect 5498 3232 5506 3296
rect 5570 3232 5586 3296
rect 5650 3232 5666 3296
rect 5730 3232 5746 3296
rect 5810 3232 5818 3296
rect 5498 3231 5818 3232
rect 14606 3296 14926 3297
rect 14606 3232 14614 3296
rect 14678 3232 14694 3296
rect 14758 3232 14774 3296
rect 14838 3232 14854 3296
rect 14918 3232 14926 3296
rect 14606 3231 14926 3232
rect 23714 3296 24034 3297
rect 23714 3232 23722 3296
rect 23786 3232 23802 3296
rect 23866 3232 23882 3296
rect 23946 3232 23962 3296
rect 24026 3232 24034 3296
rect 23714 3231 24034 3232
rect 12249 3226 12315 3229
rect 12893 3226 12959 3229
rect 12249 3224 12959 3226
rect 12249 3168 12254 3224
rect 12310 3168 12898 3224
rect 12954 3168 12959 3224
rect 12249 3166 12959 3168
rect 12249 3163 12315 3166
rect 12893 3163 12959 3166
rect 16297 3090 16363 3093
rect 20069 3090 20135 3093
rect 16297 3088 20135 3090
rect 16297 3032 16302 3088
rect 16358 3032 20074 3088
rect 20130 3032 20135 3088
rect 16297 3030 20135 3032
rect 16297 3027 16363 3030
rect 20069 3027 20135 3030
rect 12433 2954 12499 2957
rect 16665 2954 16731 2957
rect 12433 2952 16731 2954
rect 12433 2896 12438 2952
rect 12494 2896 16670 2952
rect 16726 2896 16731 2952
rect 12433 2894 16731 2896
rect 12433 2891 12499 2894
rect 16665 2891 16731 2894
rect 19333 2954 19399 2957
rect 20437 2954 20503 2957
rect 19333 2952 20503 2954
rect 19333 2896 19338 2952
rect 19394 2896 20442 2952
rect 20498 2896 20503 2952
rect 19333 2894 20503 2896
rect 19333 2891 19399 2894
rect 20437 2891 20503 2894
rect 10052 2752 10372 2753
rect 10052 2688 10060 2752
rect 10124 2688 10140 2752
rect 10204 2688 10220 2752
rect 10284 2688 10300 2752
rect 10364 2688 10372 2752
rect 10052 2687 10372 2688
rect 19160 2752 19480 2753
rect 19160 2688 19168 2752
rect 19232 2688 19248 2752
rect 19312 2688 19328 2752
rect 19392 2688 19408 2752
rect 19472 2688 19480 2752
rect 19160 2687 19480 2688
rect 9765 2412 9831 2413
rect 9765 2410 9812 2412
rect 9720 2408 9812 2410
rect 9720 2352 9770 2408
rect 9720 2350 9812 2352
rect 9765 2348 9812 2350
rect 9876 2348 9882 2412
rect 9765 2347 9831 2348
rect 5498 2208 5818 2209
rect 0 2138 800 2168
rect 5498 2144 5506 2208
rect 5570 2144 5586 2208
rect 5650 2144 5666 2208
rect 5730 2144 5746 2208
rect 5810 2144 5818 2208
rect 5498 2143 5818 2144
rect 14606 2208 14926 2209
rect 14606 2144 14614 2208
rect 14678 2144 14694 2208
rect 14758 2144 14774 2208
rect 14838 2144 14854 2208
rect 14918 2144 14926 2208
rect 14606 2143 14926 2144
rect 23714 2208 24034 2209
rect 23714 2144 23722 2208
rect 23786 2144 23802 2208
rect 23866 2144 23882 2208
rect 23946 2144 23962 2208
rect 24026 2144 24034 2208
rect 23714 2143 24034 2144
rect 2957 2138 3023 2141
rect 0 2136 3023 2138
rect 0 2080 2962 2136
rect 3018 2080 3023 2136
rect 0 2078 3023 2080
rect 0 2048 800 2078
rect 2957 2075 3023 2078
rect 26509 2138 26575 2141
rect 28780 2138 29580 2168
rect 26509 2136 29580 2138
rect 26509 2080 26514 2136
rect 26570 2080 29580 2136
rect 26509 2078 29580 2080
rect 26509 2075 26575 2078
rect 28780 2048 29580 2078
rect 0 1458 800 1488
rect 1853 1458 1919 1461
rect 0 1456 1919 1458
rect 0 1400 1858 1456
rect 1914 1400 1919 1456
rect 0 1398 1919 1400
rect 0 1368 800 1398
rect 1853 1395 1919 1398
rect 25957 1458 26023 1461
rect 28780 1458 29580 1488
rect 25957 1456 29580 1458
rect 25957 1400 25962 1456
rect 26018 1400 29580 1456
rect 25957 1398 29580 1400
rect 25957 1395 26023 1398
rect 28780 1368 29580 1398
rect 26049 778 26115 781
rect 28780 778 29580 808
rect 26049 776 29580 778
rect 26049 720 26054 776
rect 26110 720 29580 776
rect 26049 718 29580 720
rect 26049 715 26115 718
rect 28780 688 29580 718
<< via3 >>
rect 5506 29404 5570 29408
rect 5506 29348 5510 29404
rect 5510 29348 5566 29404
rect 5566 29348 5570 29404
rect 5506 29344 5570 29348
rect 5586 29404 5650 29408
rect 5586 29348 5590 29404
rect 5590 29348 5646 29404
rect 5646 29348 5650 29404
rect 5586 29344 5650 29348
rect 5666 29404 5730 29408
rect 5666 29348 5670 29404
rect 5670 29348 5726 29404
rect 5726 29348 5730 29404
rect 5666 29344 5730 29348
rect 5746 29404 5810 29408
rect 5746 29348 5750 29404
rect 5750 29348 5806 29404
rect 5806 29348 5810 29404
rect 5746 29344 5810 29348
rect 14614 29404 14678 29408
rect 14614 29348 14618 29404
rect 14618 29348 14674 29404
rect 14674 29348 14678 29404
rect 14614 29344 14678 29348
rect 14694 29404 14758 29408
rect 14694 29348 14698 29404
rect 14698 29348 14754 29404
rect 14754 29348 14758 29404
rect 14694 29344 14758 29348
rect 14774 29404 14838 29408
rect 14774 29348 14778 29404
rect 14778 29348 14834 29404
rect 14834 29348 14838 29404
rect 14774 29344 14838 29348
rect 14854 29404 14918 29408
rect 14854 29348 14858 29404
rect 14858 29348 14914 29404
rect 14914 29348 14918 29404
rect 14854 29344 14918 29348
rect 23722 29404 23786 29408
rect 23722 29348 23726 29404
rect 23726 29348 23782 29404
rect 23782 29348 23786 29404
rect 23722 29344 23786 29348
rect 23802 29404 23866 29408
rect 23802 29348 23806 29404
rect 23806 29348 23862 29404
rect 23862 29348 23866 29404
rect 23802 29344 23866 29348
rect 23882 29404 23946 29408
rect 23882 29348 23886 29404
rect 23886 29348 23942 29404
rect 23942 29348 23946 29404
rect 23882 29344 23946 29348
rect 23962 29404 24026 29408
rect 23962 29348 23966 29404
rect 23966 29348 24022 29404
rect 24022 29348 24026 29404
rect 23962 29344 24026 29348
rect 10060 28860 10124 28864
rect 10060 28804 10064 28860
rect 10064 28804 10120 28860
rect 10120 28804 10124 28860
rect 10060 28800 10124 28804
rect 10140 28860 10204 28864
rect 10140 28804 10144 28860
rect 10144 28804 10200 28860
rect 10200 28804 10204 28860
rect 10140 28800 10204 28804
rect 10220 28860 10284 28864
rect 10220 28804 10224 28860
rect 10224 28804 10280 28860
rect 10280 28804 10284 28860
rect 10220 28800 10284 28804
rect 10300 28860 10364 28864
rect 10300 28804 10304 28860
rect 10304 28804 10360 28860
rect 10360 28804 10364 28860
rect 10300 28800 10364 28804
rect 19168 28860 19232 28864
rect 19168 28804 19172 28860
rect 19172 28804 19228 28860
rect 19228 28804 19232 28860
rect 19168 28800 19232 28804
rect 19248 28860 19312 28864
rect 19248 28804 19252 28860
rect 19252 28804 19308 28860
rect 19308 28804 19312 28860
rect 19248 28800 19312 28804
rect 19328 28860 19392 28864
rect 19328 28804 19332 28860
rect 19332 28804 19388 28860
rect 19388 28804 19392 28860
rect 19328 28800 19392 28804
rect 19408 28860 19472 28864
rect 19408 28804 19412 28860
rect 19412 28804 19468 28860
rect 19468 28804 19472 28860
rect 19408 28800 19472 28804
rect 9812 28656 9876 28660
rect 9812 28600 9862 28656
rect 9862 28600 9876 28656
rect 9812 28596 9876 28600
rect 5506 28316 5570 28320
rect 5506 28260 5510 28316
rect 5510 28260 5566 28316
rect 5566 28260 5570 28316
rect 5506 28256 5570 28260
rect 5586 28316 5650 28320
rect 5586 28260 5590 28316
rect 5590 28260 5646 28316
rect 5646 28260 5650 28316
rect 5586 28256 5650 28260
rect 5666 28316 5730 28320
rect 5666 28260 5670 28316
rect 5670 28260 5726 28316
rect 5726 28260 5730 28316
rect 5666 28256 5730 28260
rect 5746 28316 5810 28320
rect 5746 28260 5750 28316
rect 5750 28260 5806 28316
rect 5806 28260 5810 28316
rect 5746 28256 5810 28260
rect 14614 28316 14678 28320
rect 14614 28260 14618 28316
rect 14618 28260 14674 28316
rect 14674 28260 14678 28316
rect 14614 28256 14678 28260
rect 14694 28316 14758 28320
rect 14694 28260 14698 28316
rect 14698 28260 14754 28316
rect 14754 28260 14758 28316
rect 14694 28256 14758 28260
rect 14774 28316 14838 28320
rect 14774 28260 14778 28316
rect 14778 28260 14834 28316
rect 14834 28260 14838 28316
rect 14774 28256 14838 28260
rect 14854 28316 14918 28320
rect 14854 28260 14858 28316
rect 14858 28260 14914 28316
rect 14914 28260 14918 28316
rect 14854 28256 14918 28260
rect 23722 28316 23786 28320
rect 23722 28260 23726 28316
rect 23726 28260 23782 28316
rect 23782 28260 23786 28316
rect 23722 28256 23786 28260
rect 23802 28316 23866 28320
rect 23802 28260 23806 28316
rect 23806 28260 23862 28316
rect 23862 28260 23866 28316
rect 23802 28256 23866 28260
rect 23882 28316 23946 28320
rect 23882 28260 23886 28316
rect 23886 28260 23942 28316
rect 23942 28260 23946 28316
rect 23882 28256 23946 28260
rect 23962 28316 24026 28320
rect 23962 28260 23966 28316
rect 23966 28260 24022 28316
rect 24022 28260 24026 28316
rect 23962 28256 24026 28260
rect 10060 27772 10124 27776
rect 10060 27716 10064 27772
rect 10064 27716 10120 27772
rect 10120 27716 10124 27772
rect 10060 27712 10124 27716
rect 10140 27772 10204 27776
rect 10140 27716 10144 27772
rect 10144 27716 10200 27772
rect 10200 27716 10204 27772
rect 10140 27712 10204 27716
rect 10220 27772 10284 27776
rect 10220 27716 10224 27772
rect 10224 27716 10280 27772
rect 10280 27716 10284 27772
rect 10220 27712 10284 27716
rect 10300 27772 10364 27776
rect 10300 27716 10304 27772
rect 10304 27716 10360 27772
rect 10360 27716 10364 27772
rect 10300 27712 10364 27716
rect 19168 27772 19232 27776
rect 19168 27716 19172 27772
rect 19172 27716 19228 27772
rect 19228 27716 19232 27772
rect 19168 27712 19232 27716
rect 19248 27772 19312 27776
rect 19248 27716 19252 27772
rect 19252 27716 19308 27772
rect 19308 27716 19312 27772
rect 19248 27712 19312 27716
rect 19328 27772 19392 27776
rect 19328 27716 19332 27772
rect 19332 27716 19388 27772
rect 19388 27716 19392 27772
rect 19328 27712 19392 27716
rect 19408 27772 19472 27776
rect 19408 27716 19412 27772
rect 19412 27716 19468 27772
rect 19468 27716 19472 27772
rect 19408 27712 19472 27716
rect 5506 27228 5570 27232
rect 5506 27172 5510 27228
rect 5510 27172 5566 27228
rect 5566 27172 5570 27228
rect 5506 27168 5570 27172
rect 5586 27228 5650 27232
rect 5586 27172 5590 27228
rect 5590 27172 5646 27228
rect 5646 27172 5650 27228
rect 5586 27168 5650 27172
rect 5666 27228 5730 27232
rect 5666 27172 5670 27228
rect 5670 27172 5726 27228
rect 5726 27172 5730 27228
rect 5666 27168 5730 27172
rect 5746 27228 5810 27232
rect 5746 27172 5750 27228
rect 5750 27172 5806 27228
rect 5806 27172 5810 27228
rect 5746 27168 5810 27172
rect 14614 27228 14678 27232
rect 14614 27172 14618 27228
rect 14618 27172 14674 27228
rect 14674 27172 14678 27228
rect 14614 27168 14678 27172
rect 14694 27228 14758 27232
rect 14694 27172 14698 27228
rect 14698 27172 14754 27228
rect 14754 27172 14758 27228
rect 14694 27168 14758 27172
rect 14774 27228 14838 27232
rect 14774 27172 14778 27228
rect 14778 27172 14834 27228
rect 14834 27172 14838 27228
rect 14774 27168 14838 27172
rect 14854 27228 14918 27232
rect 14854 27172 14858 27228
rect 14858 27172 14914 27228
rect 14914 27172 14918 27228
rect 14854 27168 14918 27172
rect 23722 27228 23786 27232
rect 23722 27172 23726 27228
rect 23726 27172 23782 27228
rect 23782 27172 23786 27228
rect 23722 27168 23786 27172
rect 23802 27228 23866 27232
rect 23802 27172 23806 27228
rect 23806 27172 23862 27228
rect 23862 27172 23866 27228
rect 23802 27168 23866 27172
rect 23882 27228 23946 27232
rect 23882 27172 23886 27228
rect 23886 27172 23942 27228
rect 23942 27172 23946 27228
rect 23882 27168 23946 27172
rect 23962 27228 24026 27232
rect 23962 27172 23966 27228
rect 23966 27172 24022 27228
rect 24022 27172 24026 27228
rect 23962 27168 24026 27172
rect 10060 26684 10124 26688
rect 10060 26628 10064 26684
rect 10064 26628 10120 26684
rect 10120 26628 10124 26684
rect 10060 26624 10124 26628
rect 10140 26684 10204 26688
rect 10140 26628 10144 26684
rect 10144 26628 10200 26684
rect 10200 26628 10204 26684
rect 10140 26624 10204 26628
rect 10220 26684 10284 26688
rect 10220 26628 10224 26684
rect 10224 26628 10280 26684
rect 10280 26628 10284 26684
rect 10220 26624 10284 26628
rect 10300 26684 10364 26688
rect 10300 26628 10304 26684
rect 10304 26628 10360 26684
rect 10360 26628 10364 26684
rect 10300 26624 10364 26628
rect 19168 26684 19232 26688
rect 19168 26628 19172 26684
rect 19172 26628 19228 26684
rect 19228 26628 19232 26684
rect 19168 26624 19232 26628
rect 19248 26684 19312 26688
rect 19248 26628 19252 26684
rect 19252 26628 19308 26684
rect 19308 26628 19312 26684
rect 19248 26624 19312 26628
rect 19328 26684 19392 26688
rect 19328 26628 19332 26684
rect 19332 26628 19388 26684
rect 19388 26628 19392 26684
rect 19328 26624 19392 26628
rect 19408 26684 19472 26688
rect 19408 26628 19412 26684
rect 19412 26628 19468 26684
rect 19468 26628 19472 26684
rect 19408 26624 19472 26628
rect 5506 26140 5570 26144
rect 5506 26084 5510 26140
rect 5510 26084 5566 26140
rect 5566 26084 5570 26140
rect 5506 26080 5570 26084
rect 5586 26140 5650 26144
rect 5586 26084 5590 26140
rect 5590 26084 5646 26140
rect 5646 26084 5650 26140
rect 5586 26080 5650 26084
rect 5666 26140 5730 26144
rect 5666 26084 5670 26140
rect 5670 26084 5726 26140
rect 5726 26084 5730 26140
rect 5666 26080 5730 26084
rect 5746 26140 5810 26144
rect 5746 26084 5750 26140
rect 5750 26084 5806 26140
rect 5806 26084 5810 26140
rect 5746 26080 5810 26084
rect 14614 26140 14678 26144
rect 14614 26084 14618 26140
rect 14618 26084 14674 26140
rect 14674 26084 14678 26140
rect 14614 26080 14678 26084
rect 14694 26140 14758 26144
rect 14694 26084 14698 26140
rect 14698 26084 14754 26140
rect 14754 26084 14758 26140
rect 14694 26080 14758 26084
rect 14774 26140 14838 26144
rect 14774 26084 14778 26140
rect 14778 26084 14834 26140
rect 14834 26084 14838 26140
rect 14774 26080 14838 26084
rect 14854 26140 14918 26144
rect 14854 26084 14858 26140
rect 14858 26084 14914 26140
rect 14914 26084 14918 26140
rect 14854 26080 14918 26084
rect 23722 26140 23786 26144
rect 23722 26084 23726 26140
rect 23726 26084 23782 26140
rect 23782 26084 23786 26140
rect 23722 26080 23786 26084
rect 23802 26140 23866 26144
rect 23802 26084 23806 26140
rect 23806 26084 23862 26140
rect 23862 26084 23866 26140
rect 23802 26080 23866 26084
rect 23882 26140 23946 26144
rect 23882 26084 23886 26140
rect 23886 26084 23942 26140
rect 23942 26084 23946 26140
rect 23882 26080 23946 26084
rect 23962 26140 24026 26144
rect 23962 26084 23966 26140
rect 23966 26084 24022 26140
rect 24022 26084 24026 26140
rect 23962 26080 24026 26084
rect 10060 25596 10124 25600
rect 10060 25540 10064 25596
rect 10064 25540 10120 25596
rect 10120 25540 10124 25596
rect 10060 25536 10124 25540
rect 10140 25596 10204 25600
rect 10140 25540 10144 25596
rect 10144 25540 10200 25596
rect 10200 25540 10204 25596
rect 10140 25536 10204 25540
rect 10220 25596 10284 25600
rect 10220 25540 10224 25596
rect 10224 25540 10280 25596
rect 10280 25540 10284 25596
rect 10220 25536 10284 25540
rect 10300 25596 10364 25600
rect 10300 25540 10304 25596
rect 10304 25540 10360 25596
rect 10360 25540 10364 25596
rect 10300 25536 10364 25540
rect 19168 25596 19232 25600
rect 19168 25540 19172 25596
rect 19172 25540 19228 25596
rect 19228 25540 19232 25596
rect 19168 25536 19232 25540
rect 19248 25596 19312 25600
rect 19248 25540 19252 25596
rect 19252 25540 19308 25596
rect 19308 25540 19312 25596
rect 19248 25536 19312 25540
rect 19328 25596 19392 25600
rect 19328 25540 19332 25596
rect 19332 25540 19388 25596
rect 19388 25540 19392 25596
rect 19328 25536 19392 25540
rect 19408 25596 19472 25600
rect 19408 25540 19412 25596
rect 19412 25540 19468 25596
rect 19468 25540 19472 25596
rect 19408 25536 19472 25540
rect 5506 25052 5570 25056
rect 5506 24996 5510 25052
rect 5510 24996 5566 25052
rect 5566 24996 5570 25052
rect 5506 24992 5570 24996
rect 5586 25052 5650 25056
rect 5586 24996 5590 25052
rect 5590 24996 5646 25052
rect 5646 24996 5650 25052
rect 5586 24992 5650 24996
rect 5666 25052 5730 25056
rect 5666 24996 5670 25052
rect 5670 24996 5726 25052
rect 5726 24996 5730 25052
rect 5666 24992 5730 24996
rect 5746 25052 5810 25056
rect 5746 24996 5750 25052
rect 5750 24996 5806 25052
rect 5806 24996 5810 25052
rect 5746 24992 5810 24996
rect 14614 25052 14678 25056
rect 14614 24996 14618 25052
rect 14618 24996 14674 25052
rect 14674 24996 14678 25052
rect 14614 24992 14678 24996
rect 14694 25052 14758 25056
rect 14694 24996 14698 25052
rect 14698 24996 14754 25052
rect 14754 24996 14758 25052
rect 14694 24992 14758 24996
rect 14774 25052 14838 25056
rect 14774 24996 14778 25052
rect 14778 24996 14834 25052
rect 14834 24996 14838 25052
rect 14774 24992 14838 24996
rect 14854 25052 14918 25056
rect 14854 24996 14858 25052
rect 14858 24996 14914 25052
rect 14914 24996 14918 25052
rect 14854 24992 14918 24996
rect 23722 25052 23786 25056
rect 23722 24996 23726 25052
rect 23726 24996 23782 25052
rect 23782 24996 23786 25052
rect 23722 24992 23786 24996
rect 23802 25052 23866 25056
rect 23802 24996 23806 25052
rect 23806 24996 23862 25052
rect 23862 24996 23866 25052
rect 23802 24992 23866 24996
rect 23882 25052 23946 25056
rect 23882 24996 23886 25052
rect 23886 24996 23942 25052
rect 23942 24996 23946 25052
rect 23882 24992 23946 24996
rect 23962 25052 24026 25056
rect 23962 24996 23966 25052
rect 23966 24996 24022 25052
rect 24022 24996 24026 25052
rect 23962 24992 24026 24996
rect 10060 24508 10124 24512
rect 10060 24452 10064 24508
rect 10064 24452 10120 24508
rect 10120 24452 10124 24508
rect 10060 24448 10124 24452
rect 10140 24508 10204 24512
rect 10140 24452 10144 24508
rect 10144 24452 10200 24508
rect 10200 24452 10204 24508
rect 10140 24448 10204 24452
rect 10220 24508 10284 24512
rect 10220 24452 10224 24508
rect 10224 24452 10280 24508
rect 10280 24452 10284 24508
rect 10220 24448 10284 24452
rect 10300 24508 10364 24512
rect 10300 24452 10304 24508
rect 10304 24452 10360 24508
rect 10360 24452 10364 24508
rect 10300 24448 10364 24452
rect 19168 24508 19232 24512
rect 19168 24452 19172 24508
rect 19172 24452 19228 24508
rect 19228 24452 19232 24508
rect 19168 24448 19232 24452
rect 19248 24508 19312 24512
rect 19248 24452 19252 24508
rect 19252 24452 19308 24508
rect 19308 24452 19312 24508
rect 19248 24448 19312 24452
rect 19328 24508 19392 24512
rect 19328 24452 19332 24508
rect 19332 24452 19388 24508
rect 19388 24452 19392 24508
rect 19328 24448 19392 24452
rect 19408 24508 19472 24512
rect 19408 24452 19412 24508
rect 19412 24452 19468 24508
rect 19468 24452 19472 24508
rect 19408 24448 19472 24452
rect 9812 24168 9876 24172
rect 9812 24112 9862 24168
rect 9862 24112 9876 24168
rect 9812 24108 9876 24112
rect 5506 23964 5570 23968
rect 5506 23908 5510 23964
rect 5510 23908 5566 23964
rect 5566 23908 5570 23964
rect 5506 23904 5570 23908
rect 5586 23964 5650 23968
rect 5586 23908 5590 23964
rect 5590 23908 5646 23964
rect 5646 23908 5650 23964
rect 5586 23904 5650 23908
rect 5666 23964 5730 23968
rect 5666 23908 5670 23964
rect 5670 23908 5726 23964
rect 5726 23908 5730 23964
rect 5666 23904 5730 23908
rect 5746 23964 5810 23968
rect 5746 23908 5750 23964
rect 5750 23908 5806 23964
rect 5806 23908 5810 23964
rect 5746 23904 5810 23908
rect 14614 23964 14678 23968
rect 14614 23908 14618 23964
rect 14618 23908 14674 23964
rect 14674 23908 14678 23964
rect 14614 23904 14678 23908
rect 14694 23964 14758 23968
rect 14694 23908 14698 23964
rect 14698 23908 14754 23964
rect 14754 23908 14758 23964
rect 14694 23904 14758 23908
rect 14774 23964 14838 23968
rect 14774 23908 14778 23964
rect 14778 23908 14834 23964
rect 14834 23908 14838 23964
rect 14774 23904 14838 23908
rect 14854 23964 14918 23968
rect 14854 23908 14858 23964
rect 14858 23908 14914 23964
rect 14914 23908 14918 23964
rect 14854 23904 14918 23908
rect 23722 23964 23786 23968
rect 23722 23908 23726 23964
rect 23726 23908 23782 23964
rect 23782 23908 23786 23964
rect 23722 23904 23786 23908
rect 23802 23964 23866 23968
rect 23802 23908 23806 23964
rect 23806 23908 23862 23964
rect 23862 23908 23866 23964
rect 23802 23904 23866 23908
rect 23882 23964 23946 23968
rect 23882 23908 23886 23964
rect 23886 23908 23942 23964
rect 23942 23908 23946 23964
rect 23882 23904 23946 23908
rect 23962 23964 24026 23968
rect 23962 23908 23966 23964
rect 23966 23908 24022 23964
rect 24022 23908 24026 23964
rect 23962 23904 24026 23908
rect 26372 23488 26436 23492
rect 26372 23432 26386 23488
rect 26386 23432 26436 23488
rect 26372 23428 26436 23432
rect 10060 23420 10124 23424
rect 10060 23364 10064 23420
rect 10064 23364 10120 23420
rect 10120 23364 10124 23420
rect 10060 23360 10124 23364
rect 10140 23420 10204 23424
rect 10140 23364 10144 23420
rect 10144 23364 10200 23420
rect 10200 23364 10204 23420
rect 10140 23360 10204 23364
rect 10220 23420 10284 23424
rect 10220 23364 10224 23420
rect 10224 23364 10280 23420
rect 10280 23364 10284 23420
rect 10220 23360 10284 23364
rect 10300 23420 10364 23424
rect 10300 23364 10304 23420
rect 10304 23364 10360 23420
rect 10360 23364 10364 23420
rect 10300 23360 10364 23364
rect 19168 23420 19232 23424
rect 19168 23364 19172 23420
rect 19172 23364 19228 23420
rect 19228 23364 19232 23420
rect 19168 23360 19232 23364
rect 19248 23420 19312 23424
rect 19248 23364 19252 23420
rect 19252 23364 19308 23420
rect 19308 23364 19312 23420
rect 19248 23360 19312 23364
rect 19328 23420 19392 23424
rect 19328 23364 19332 23420
rect 19332 23364 19388 23420
rect 19388 23364 19392 23420
rect 19328 23360 19392 23364
rect 19408 23420 19472 23424
rect 19408 23364 19412 23420
rect 19412 23364 19468 23420
rect 19468 23364 19472 23420
rect 19408 23360 19472 23364
rect 5506 22876 5570 22880
rect 5506 22820 5510 22876
rect 5510 22820 5566 22876
rect 5566 22820 5570 22876
rect 5506 22816 5570 22820
rect 5586 22876 5650 22880
rect 5586 22820 5590 22876
rect 5590 22820 5646 22876
rect 5646 22820 5650 22876
rect 5586 22816 5650 22820
rect 5666 22876 5730 22880
rect 5666 22820 5670 22876
rect 5670 22820 5726 22876
rect 5726 22820 5730 22876
rect 5666 22816 5730 22820
rect 5746 22876 5810 22880
rect 5746 22820 5750 22876
rect 5750 22820 5806 22876
rect 5806 22820 5810 22876
rect 5746 22816 5810 22820
rect 14614 22876 14678 22880
rect 14614 22820 14618 22876
rect 14618 22820 14674 22876
rect 14674 22820 14678 22876
rect 14614 22816 14678 22820
rect 14694 22876 14758 22880
rect 14694 22820 14698 22876
rect 14698 22820 14754 22876
rect 14754 22820 14758 22876
rect 14694 22816 14758 22820
rect 14774 22876 14838 22880
rect 14774 22820 14778 22876
rect 14778 22820 14834 22876
rect 14834 22820 14838 22876
rect 14774 22816 14838 22820
rect 14854 22876 14918 22880
rect 14854 22820 14858 22876
rect 14858 22820 14914 22876
rect 14914 22820 14918 22876
rect 14854 22816 14918 22820
rect 23722 22876 23786 22880
rect 23722 22820 23726 22876
rect 23726 22820 23782 22876
rect 23782 22820 23786 22876
rect 23722 22816 23786 22820
rect 23802 22876 23866 22880
rect 23802 22820 23806 22876
rect 23806 22820 23862 22876
rect 23862 22820 23866 22876
rect 23802 22816 23866 22820
rect 23882 22876 23946 22880
rect 23882 22820 23886 22876
rect 23886 22820 23942 22876
rect 23942 22820 23946 22876
rect 23882 22816 23946 22820
rect 23962 22876 24026 22880
rect 23962 22820 23966 22876
rect 23966 22820 24022 22876
rect 24022 22820 24026 22876
rect 23962 22816 24026 22820
rect 10060 22332 10124 22336
rect 10060 22276 10064 22332
rect 10064 22276 10120 22332
rect 10120 22276 10124 22332
rect 10060 22272 10124 22276
rect 10140 22332 10204 22336
rect 10140 22276 10144 22332
rect 10144 22276 10200 22332
rect 10200 22276 10204 22332
rect 10140 22272 10204 22276
rect 10220 22332 10284 22336
rect 10220 22276 10224 22332
rect 10224 22276 10280 22332
rect 10280 22276 10284 22332
rect 10220 22272 10284 22276
rect 10300 22332 10364 22336
rect 10300 22276 10304 22332
rect 10304 22276 10360 22332
rect 10360 22276 10364 22332
rect 10300 22272 10364 22276
rect 19168 22332 19232 22336
rect 19168 22276 19172 22332
rect 19172 22276 19228 22332
rect 19228 22276 19232 22332
rect 19168 22272 19232 22276
rect 19248 22332 19312 22336
rect 19248 22276 19252 22332
rect 19252 22276 19308 22332
rect 19308 22276 19312 22332
rect 19248 22272 19312 22276
rect 19328 22332 19392 22336
rect 19328 22276 19332 22332
rect 19332 22276 19388 22332
rect 19388 22276 19392 22332
rect 19328 22272 19392 22276
rect 19408 22332 19472 22336
rect 19408 22276 19412 22332
rect 19412 22276 19468 22332
rect 19468 22276 19472 22332
rect 19408 22272 19472 22276
rect 5506 21788 5570 21792
rect 5506 21732 5510 21788
rect 5510 21732 5566 21788
rect 5566 21732 5570 21788
rect 5506 21728 5570 21732
rect 5586 21788 5650 21792
rect 5586 21732 5590 21788
rect 5590 21732 5646 21788
rect 5646 21732 5650 21788
rect 5586 21728 5650 21732
rect 5666 21788 5730 21792
rect 5666 21732 5670 21788
rect 5670 21732 5726 21788
rect 5726 21732 5730 21788
rect 5666 21728 5730 21732
rect 5746 21788 5810 21792
rect 5746 21732 5750 21788
rect 5750 21732 5806 21788
rect 5806 21732 5810 21788
rect 5746 21728 5810 21732
rect 14614 21788 14678 21792
rect 14614 21732 14618 21788
rect 14618 21732 14674 21788
rect 14674 21732 14678 21788
rect 14614 21728 14678 21732
rect 14694 21788 14758 21792
rect 14694 21732 14698 21788
rect 14698 21732 14754 21788
rect 14754 21732 14758 21788
rect 14694 21728 14758 21732
rect 14774 21788 14838 21792
rect 14774 21732 14778 21788
rect 14778 21732 14834 21788
rect 14834 21732 14838 21788
rect 14774 21728 14838 21732
rect 14854 21788 14918 21792
rect 14854 21732 14858 21788
rect 14858 21732 14914 21788
rect 14914 21732 14918 21788
rect 14854 21728 14918 21732
rect 23722 21788 23786 21792
rect 23722 21732 23726 21788
rect 23726 21732 23782 21788
rect 23782 21732 23786 21788
rect 23722 21728 23786 21732
rect 23802 21788 23866 21792
rect 23802 21732 23806 21788
rect 23806 21732 23862 21788
rect 23862 21732 23866 21788
rect 23802 21728 23866 21732
rect 23882 21788 23946 21792
rect 23882 21732 23886 21788
rect 23886 21732 23942 21788
rect 23942 21732 23946 21788
rect 23882 21728 23946 21732
rect 23962 21788 24026 21792
rect 23962 21732 23966 21788
rect 23966 21732 24022 21788
rect 24022 21732 24026 21788
rect 23962 21728 24026 21732
rect 10060 21244 10124 21248
rect 10060 21188 10064 21244
rect 10064 21188 10120 21244
rect 10120 21188 10124 21244
rect 10060 21184 10124 21188
rect 10140 21244 10204 21248
rect 10140 21188 10144 21244
rect 10144 21188 10200 21244
rect 10200 21188 10204 21244
rect 10140 21184 10204 21188
rect 10220 21244 10284 21248
rect 10220 21188 10224 21244
rect 10224 21188 10280 21244
rect 10280 21188 10284 21244
rect 10220 21184 10284 21188
rect 10300 21244 10364 21248
rect 10300 21188 10304 21244
rect 10304 21188 10360 21244
rect 10360 21188 10364 21244
rect 10300 21184 10364 21188
rect 19168 21244 19232 21248
rect 19168 21188 19172 21244
rect 19172 21188 19228 21244
rect 19228 21188 19232 21244
rect 19168 21184 19232 21188
rect 19248 21244 19312 21248
rect 19248 21188 19252 21244
rect 19252 21188 19308 21244
rect 19308 21188 19312 21244
rect 19248 21184 19312 21188
rect 19328 21244 19392 21248
rect 19328 21188 19332 21244
rect 19332 21188 19388 21244
rect 19388 21188 19392 21244
rect 19328 21184 19392 21188
rect 19408 21244 19472 21248
rect 19408 21188 19412 21244
rect 19412 21188 19468 21244
rect 19468 21188 19472 21244
rect 19408 21184 19472 21188
rect 5506 20700 5570 20704
rect 5506 20644 5510 20700
rect 5510 20644 5566 20700
rect 5566 20644 5570 20700
rect 5506 20640 5570 20644
rect 5586 20700 5650 20704
rect 5586 20644 5590 20700
rect 5590 20644 5646 20700
rect 5646 20644 5650 20700
rect 5586 20640 5650 20644
rect 5666 20700 5730 20704
rect 5666 20644 5670 20700
rect 5670 20644 5726 20700
rect 5726 20644 5730 20700
rect 5666 20640 5730 20644
rect 5746 20700 5810 20704
rect 5746 20644 5750 20700
rect 5750 20644 5806 20700
rect 5806 20644 5810 20700
rect 5746 20640 5810 20644
rect 14614 20700 14678 20704
rect 14614 20644 14618 20700
rect 14618 20644 14674 20700
rect 14674 20644 14678 20700
rect 14614 20640 14678 20644
rect 14694 20700 14758 20704
rect 14694 20644 14698 20700
rect 14698 20644 14754 20700
rect 14754 20644 14758 20700
rect 14694 20640 14758 20644
rect 14774 20700 14838 20704
rect 14774 20644 14778 20700
rect 14778 20644 14834 20700
rect 14834 20644 14838 20700
rect 14774 20640 14838 20644
rect 14854 20700 14918 20704
rect 14854 20644 14858 20700
rect 14858 20644 14914 20700
rect 14914 20644 14918 20700
rect 14854 20640 14918 20644
rect 23722 20700 23786 20704
rect 23722 20644 23726 20700
rect 23726 20644 23782 20700
rect 23782 20644 23786 20700
rect 23722 20640 23786 20644
rect 23802 20700 23866 20704
rect 23802 20644 23806 20700
rect 23806 20644 23862 20700
rect 23862 20644 23866 20700
rect 23802 20640 23866 20644
rect 23882 20700 23946 20704
rect 23882 20644 23886 20700
rect 23886 20644 23942 20700
rect 23942 20644 23946 20700
rect 23882 20640 23946 20644
rect 23962 20700 24026 20704
rect 23962 20644 23966 20700
rect 23966 20644 24022 20700
rect 24022 20644 24026 20700
rect 23962 20640 24026 20644
rect 10060 20156 10124 20160
rect 10060 20100 10064 20156
rect 10064 20100 10120 20156
rect 10120 20100 10124 20156
rect 10060 20096 10124 20100
rect 10140 20156 10204 20160
rect 10140 20100 10144 20156
rect 10144 20100 10200 20156
rect 10200 20100 10204 20156
rect 10140 20096 10204 20100
rect 10220 20156 10284 20160
rect 10220 20100 10224 20156
rect 10224 20100 10280 20156
rect 10280 20100 10284 20156
rect 10220 20096 10284 20100
rect 10300 20156 10364 20160
rect 10300 20100 10304 20156
rect 10304 20100 10360 20156
rect 10360 20100 10364 20156
rect 10300 20096 10364 20100
rect 19168 20156 19232 20160
rect 19168 20100 19172 20156
rect 19172 20100 19228 20156
rect 19228 20100 19232 20156
rect 19168 20096 19232 20100
rect 19248 20156 19312 20160
rect 19248 20100 19252 20156
rect 19252 20100 19308 20156
rect 19308 20100 19312 20156
rect 19248 20096 19312 20100
rect 19328 20156 19392 20160
rect 19328 20100 19332 20156
rect 19332 20100 19388 20156
rect 19388 20100 19392 20156
rect 19328 20096 19392 20100
rect 19408 20156 19472 20160
rect 19408 20100 19412 20156
rect 19412 20100 19468 20156
rect 19468 20100 19472 20156
rect 19408 20096 19472 20100
rect 5506 19612 5570 19616
rect 5506 19556 5510 19612
rect 5510 19556 5566 19612
rect 5566 19556 5570 19612
rect 5506 19552 5570 19556
rect 5586 19612 5650 19616
rect 5586 19556 5590 19612
rect 5590 19556 5646 19612
rect 5646 19556 5650 19612
rect 5586 19552 5650 19556
rect 5666 19612 5730 19616
rect 5666 19556 5670 19612
rect 5670 19556 5726 19612
rect 5726 19556 5730 19612
rect 5666 19552 5730 19556
rect 5746 19612 5810 19616
rect 5746 19556 5750 19612
rect 5750 19556 5806 19612
rect 5806 19556 5810 19612
rect 5746 19552 5810 19556
rect 14614 19612 14678 19616
rect 14614 19556 14618 19612
rect 14618 19556 14674 19612
rect 14674 19556 14678 19612
rect 14614 19552 14678 19556
rect 14694 19612 14758 19616
rect 14694 19556 14698 19612
rect 14698 19556 14754 19612
rect 14754 19556 14758 19612
rect 14694 19552 14758 19556
rect 14774 19612 14838 19616
rect 14774 19556 14778 19612
rect 14778 19556 14834 19612
rect 14834 19556 14838 19612
rect 14774 19552 14838 19556
rect 14854 19612 14918 19616
rect 14854 19556 14858 19612
rect 14858 19556 14914 19612
rect 14914 19556 14918 19612
rect 14854 19552 14918 19556
rect 23722 19612 23786 19616
rect 23722 19556 23726 19612
rect 23726 19556 23782 19612
rect 23782 19556 23786 19612
rect 23722 19552 23786 19556
rect 23802 19612 23866 19616
rect 23802 19556 23806 19612
rect 23806 19556 23862 19612
rect 23862 19556 23866 19612
rect 23802 19552 23866 19556
rect 23882 19612 23946 19616
rect 23882 19556 23886 19612
rect 23886 19556 23942 19612
rect 23942 19556 23946 19612
rect 23882 19552 23946 19556
rect 23962 19612 24026 19616
rect 23962 19556 23966 19612
rect 23966 19556 24022 19612
rect 24022 19556 24026 19612
rect 23962 19552 24026 19556
rect 9812 19212 9876 19276
rect 10060 19068 10124 19072
rect 10060 19012 10064 19068
rect 10064 19012 10120 19068
rect 10120 19012 10124 19068
rect 10060 19008 10124 19012
rect 10140 19068 10204 19072
rect 10140 19012 10144 19068
rect 10144 19012 10200 19068
rect 10200 19012 10204 19068
rect 10140 19008 10204 19012
rect 10220 19068 10284 19072
rect 10220 19012 10224 19068
rect 10224 19012 10280 19068
rect 10280 19012 10284 19068
rect 10220 19008 10284 19012
rect 10300 19068 10364 19072
rect 10300 19012 10304 19068
rect 10304 19012 10360 19068
rect 10360 19012 10364 19068
rect 10300 19008 10364 19012
rect 19168 19068 19232 19072
rect 19168 19012 19172 19068
rect 19172 19012 19228 19068
rect 19228 19012 19232 19068
rect 19168 19008 19232 19012
rect 19248 19068 19312 19072
rect 19248 19012 19252 19068
rect 19252 19012 19308 19068
rect 19308 19012 19312 19068
rect 19248 19008 19312 19012
rect 19328 19068 19392 19072
rect 19328 19012 19332 19068
rect 19332 19012 19388 19068
rect 19388 19012 19392 19068
rect 19328 19008 19392 19012
rect 19408 19068 19472 19072
rect 19408 19012 19412 19068
rect 19412 19012 19468 19068
rect 19468 19012 19472 19068
rect 19408 19008 19472 19012
rect 5506 18524 5570 18528
rect 5506 18468 5510 18524
rect 5510 18468 5566 18524
rect 5566 18468 5570 18524
rect 5506 18464 5570 18468
rect 5586 18524 5650 18528
rect 5586 18468 5590 18524
rect 5590 18468 5646 18524
rect 5646 18468 5650 18524
rect 5586 18464 5650 18468
rect 5666 18524 5730 18528
rect 5666 18468 5670 18524
rect 5670 18468 5726 18524
rect 5726 18468 5730 18524
rect 5666 18464 5730 18468
rect 5746 18524 5810 18528
rect 5746 18468 5750 18524
rect 5750 18468 5806 18524
rect 5806 18468 5810 18524
rect 5746 18464 5810 18468
rect 14614 18524 14678 18528
rect 14614 18468 14618 18524
rect 14618 18468 14674 18524
rect 14674 18468 14678 18524
rect 14614 18464 14678 18468
rect 14694 18524 14758 18528
rect 14694 18468 14698 18524
rect 14698 18468 14754 18524
rect 14754 18468 14758 18524
rect 14694 18464 14758 18468
rect 14774 18524 14838 18528
rect 14774 18468 14778 18524
rect 14778 18468 14834 18524
rect 14834 18468 14838 18524
rect 14774 18464 14838 18468
rect 14854 18524 14918 18528
rect 14854 18468 14858 18524
rect 14858 18468 14914 18524
rect 14914 18468 14918 18524
rect 14854 18464 14918 18468
rect 23722 18524 23786 18528
rect 23722 18468 23726 18524
rect 23726 18468 23782 18524
rect 23782 18468 23786 18524
rect 23722 18464 23786 18468
rect 23802 18524 23866 18528
rect 23802 18468 23806 18524
rect 23806 18468 23862 18524
rect 23862 18468 23866 18524
rect 23802 18464 23866 18468
rect 23882 18524 23946 18528
rect 23882 18468 23886 18524
rect 23886 18468 23942 18524
rect 23942 18468 23946 18524
rect 23882 18464 23946 18468
rect 23962 18524 24026 18528
rect 23962 18468 23966 18524
rect 23966 18468 24022 18524
rect 24022 18468 24026 18524
rect 23962 18464 24026 18468
rect 10060 17980 10124 17984
rect 10060 17924 10064 17980
rect 10064 17924 10120 17980
rect 10120 17924 10124 17980
rect 10060 17920 10124 17924
rect 10140 17980 10204 17984
rect 10140 17924 10144 17980
rect 10144 17924 10200 17980
rect 10200 17924 10204 17980
rect 10140 17920 10204 17924
rect 10220 17980 10284 17984
rect 10220 17924 10224 17980
rect 10224 17924 10280 17980
rect 10280 17924 10284 17980
rect 10220 17920 10284 17924
rect 10300 17980 10364 17984
rect 10300 17924 10304 17980
rect 10304 17924 10360 17980
rect 10360 17924 10364 17980
rect 10300 17920 10364 17924
rect 19168 17980 19232 17984
rect 19168 17924 19172 17980
rect 19172 17924 19228 17980
rect 19228 17924 19232 17980
rect 19168 17920 19232 17924
rect 19248 17980 19312 17984
rect 19248 17924 19252 17980
rect 19252 17924 19308 17980
rect 19308 17924 19312 17980
rect 19248 17920 19312 17924
rect 19328 17980 19392 17984
rect 19328 17924 19332 17980
rect 19332 17924 19388 17980
rect 19388 17924 19392 17980
rect 19328 17920 19392 17924
rect 19408 17980 19472 17984
rect 19408 17924 19412 17980
rect 19412 17924 19468 17980
rect 19468 17924 19472 17980
rect 19408 17920 19472 17924
rect 5506 17436 5570 17440
rect 5506 17380 5510 17436
rect 5510 17380 5566 17436
rect 5566 17380 5570 17436
rect 5506 17376 5570 17380
rect 5586 17436 5650 17440
rect 5586 17380 5590 17436
rect 5590 17380 5646 17436
rect 5646 17380 5650 17436
rect 5586 17376 5650 17380
rect 5666 17436 5730 17440
rect 5666 17380 5670 17436
rect 5670 17380 5726 17436
rect 5726 17380 5730 17436
rect 5666 17376 5730 17380
rect 5746 17436 5810 17440
rect 5746 17380 5750 17436
rect 5750 17380 5806 17436
rect 5806 17380 5810 17436
rect 5746 17376 5810 17380
rect 14614 17436 14678 17440
rect 14614 17380 14618 17436
rect 14618 17380 14674 17436
rect 14674 17380 14678 17436
rect 14614 17376 14678 17380
rect 14694 17436 14758 17440
rect 14694 17380 14698 17436
rect 14698 17380 14754 17436
rect 14754 17380 14758 17436
rect 14694 17376 14758 17380
rect 14774 17436 14838 17440
rect 14774 17380 14778 17436
rect 14778 17380 14834 17436
rect 14834 17380 14838 17436
rect 14774 17376 14838 17380
rect 14854 17436 14918 17440
rect 14854 17380 14858 17436
rect 14858 17380 14914 17436
rect 14914 17380 14918 17436
rect 14854 17376 14918 17380
rect 23722 17436 23786 17440
rect 23722 17380 23726 17436
rect 23726 17380 23782 17436
rect 23782 17380 23786 17436
rect 23722 17376 23786 17380
rect 23802 17436 23866 17440
rect 23802 17380 23806 17436
rect 23806 17380 23862 17436
rect 23862 17380 23866 17436
rect 23802 17376 23866 17380
rect 23882 17436 23946 17440
rect 23882 17380 23886 17436
rect 23886 17380 23942 17436
rect 23942 17380 23946 17436
rect 23882 17376 23946 17380
rect 23962 17436 24026 17440
rect 23962 17380 23966 17436
rect 23966 17380 24022 17436
rect 24022 17380 24026 17436
rect 23962 17376 24026 17380
rect 9812 17368 9876 17372
rect 9812 17312 9862 17368
rect 9862 17312 9876 17368
rect 9812 17308 9876 17312
rect 10060 16892 10124 16896
rect 10060 16836 10064 16892
rect 10064 16836 10120 16892
rect 10120 16836 10124 16892
rect 10060 16832 10124 16836
rect 10140 16892 10204 16896
rect 10140 16836 10144 16892
rect 10144 16836 10200 16892
rect 10200 16836 10204 16892
rect 10140 16832 10204 16836
rect 10220 16892 10284 16896
rect 10220 16836 10224 16892
rect 10224 16836 10280 16892
rect 10280 16836 10284 16892
rect 10220 16832 10284 16836
rect 10300 16892 10364 16896
rect 10300 16836 10304 16892
rect 10304 16836 10360 16892
rect 10360 16836 10364 16892
rect 10300 16832 10364 16836
rect 19168 16892 19232 16896
rect 19168 16836 19172 16892
rect 19172 16836 19228 16892
rect 19228 16836 19232 16892
rect 19168 16832 19232 16836
rect 19248 16892 19312 16896
rect 19248 16836 19252 16892
rect 19252 16836 19308 16892
rect 19308 16836 19312 16892
rect 19248 16832 19312 16836
rect 19328 16892 19392 16896
rect 19328 16836 19332 16892
rect 19332 16836 19388 16892
rect 19388 16836 19392 16892
rect 19328 16832 19392 16836
rect 19408 16892 19472 16896
rect 19408 16836 19412 16892
rect 19412 16836 19468 16892
rect 19468 16836 19472 16892
rect 19408 16832 19472 16836
rect 5506 16348 5570 16352
rect 5506 16292 5510 16348
rect 5510 16292 5566 16348
rect 5566 16292 5570 16348
rect 5506 16288 5570 16292
rect 5586 16348 5650 16352
rect 5586 16292 5590 16348
rect 5590 16292 5646 16348
rect 5646 16292 5650 16348
rect 5586 16288 5650 16292
rect 5666 16348 5730 16352
rect 5666 16292 5670 16348
rect 5670 16292 5726 16348
rect 5726 16292 5730 16348
rect 5666 16288 5730 16292
rect 5746 16348 5810 16352
rect 5746 16292 5750 16348
rect 5750 16292 5806 16348
rect 5806 16292 5810 16348
rect 5746 16288 5810 16292
rect 14614 16348 14678 16352
rect 14614 16292 14618 16348
rect 14618 16292 14674 16348
rect 14674 16292 14678 16348
rect 14614 16288 14678 16292
rect 14694 16348 14758 16352
rect 14694 16292 14698 16348
rect 14698 16292 14754 16348
rect 14754 16292 14758 16348
rect 14694 16288 14758 16292
rect 14774 16348 14838 16352
rect 14774 16292 14778 16348
rect 14778 16292 14834 16348
rect 14834 16292 14838 16348
rect 14774 16288 14838 16292
rect 14854 16348 14918 16352
rect 14854 16292 14858 16348
rect 14858 16292 14914 16348
rect 14914 16292 14918 16348
rect 14854 16288 14918 16292
rect 23722 16348 23786 16352
rect 23722 16292 23726 16348
rect 23726 16292 23782 16348
rect 23782 16292 23786 16348
rect 23722 16288 23786 16292
rect 23802 16348 23866 16352
rect 23802 16292 23806 16348
rect 23806 16292 23862 16348
rect 23862 16292 23866 16348
rect 23802 16288 23866 16292
rect 23882 16348 23946 16352
rect 23882 16292 23886 16348
rect 23886 16292 23942 16348
rect 23942 16292 23946 16348
rect 23882 16288 23946 16292
rect 23962 16348 24026 16352
rect 23962 16292 23966 16348
rect 23966 16292 24022 16348
rect 24022 16292 24026 16348
rect 23962 16288 24026 16292
rect 10916 16084 10980 16148
rect 10060 15804 10124 15808
rect 10060 15748 10064 15804
rect 10064 15748 10120 15804
rect 10120 15748 10124 15804
rect 10060 15744 10124 15748
rect 10140 15804 10204 15808
rect 10140 15748 10144 15804
rect 10144 15748 10200 15804
rect 10200 15748 10204 15804
rect 10140 15744 10204 15748
rect 10220 15804 10284 15808
rect 10220 15748 10224 15804
rect 10224 15748 10280 15804
rect 10280 15748 10284 15804
rect 10220 15744 10284 15748
rect 10300 15804 10364 15808
rect 10300 15748 10304 15804
rect 10304 15748 10360 15804
rect 10360 15748 10364 15804
rect 10300 15744 10364 15748
rect 19168 15804 19232 15808
rect 19168 15748 19172 15804
rect 19172 15748 19228 15804
rect 19228 15748 19232 15804
rect 19168 15744 19232 15748
rect 19248 15804 19312 15808
rect 19248 15748 19252 15804
rect 19252 15748 19308 15804
rect 19308 15748 19312 15804
rect 19248 15744 19312 15748
rect 19328 15804 19392 15808
rect 19328 15748 19332 15804
rect 19332 15748 19388 15804
rect 19388 15748 19392 15804
rect 19328 15744 19392 15748
rect 19408 15804 19472 15808
rect 19408 15748 19412 15804
rect 19412 15748 19468 15804
rect 19468 15748 19472 15804
rect 19408 15744 19472 15748
rect 5506 15260 5570 15264
rect 5506 15204 5510 15260
rect 5510 15204 5566 15260
rect 5566 15204 5570 15260
rect 5506 15200 5570 15204
rect 5586 15260 5650 15264
rect 5586 15204 5590 15260
rect 5590 15204 5646 15260
rect 5646 15204 5650 15260
rect 5586 15200 5650 15204
rect 5666 15260 5730 15264
rect 5666 15204 5670 15260
rect 5670 15204 5726 15260
rect 5726 15204 5730 15260
rect 5666 15200 5730 15204
rect 5746 15260 5810 15264
rect 5746 15204 5750 15260
rect 5750 15204 5806 15260
rect 5806 15204 5810 15260
rect 5746 15200 5810 15204
rect 14614 15260 14678 15264
rect 14614 15204 14618 15260
rect 14618 15204 14674 15260
rect 14674 15204 14678 15260
rect 14614 15200 14678 15204
rect 14694 15260 14758 15264
rect 14694 15204 14698 15260
rect 14698 15204 14754 15260
rect 14754 15204 14758 15260
rect 14694 15200 14758 15204
rect 14774 15260 14838 15264
rect 14774 15204 14778 15260
rect 14778 15204 14834 15260
rect 14834 15204 14838 15260
rect 14774 15200 14838 15204
rect 14854 15260 14918 15264
rect 14854 15204 14858 15260
rect 14858 15204 14914 15260
rect 14914 15204 14918 15260
rect 14854 15200 14918 15204
rect 23722 15260 23786 15264
rect 23722 15204 23726 15260
rect 23726 15204 23782 15260
rect 23782 15204 23786 15260
rect 23722 15200 23786 15204
rect 23802 15260 23866 15264
rect 23802 15204 23806 15260
rect 23806 15204 23862 15260
rect 23862 15204 23866 15260
rect 23802 15200 23866 15204
rect 23882 15260 23946 15264
rect 23882 15204 23886 15260
rect 23886 15204 23942 15260
rect 23942 15204 23946 15260
rect 23882 15200 23946 15204
rect 23962 15260 24026 15264
rect 23962 15204 23966 15260
rect 23966 15204 24022 15260
rect 24022 15204 24026 15260
rect 23962 15200 24026 15204
rect 10060 14716 10124 14720
rect 10060 14660 10064 14716
rect 10064 14660 10120 14716
rect 10120 14660 10124 14716
rect 10060 14656 10124 14660
rect 10140 14716 10204 14720
rect 10140 14660 10144 14716
rect 10144 14660 10200 14716
rect 10200 14660 10204 14716
rect 10140 14656 10204 14660
rect 10220 14716 10284 14720
rect 10220 14660 10224 14716
rect 10224 14660 10280 14716
rect 10280 14660 10284 14716
rect 10220 14656 10284 14660
rect 10300 14716 10364 14720
rect 10300 14660 10304 14716
rect 10304 14660 10360 14716
rect 10360 14660 10364 14716
rect 10300 14656 10364 14660
rect 19168 14716 19232 14720
rect 19168 14660 19172 14716
rect 19172 14660 19228 14716
rect 19228 14660 19232 14716
rect 19168 14656 19232 14660
rect 19248 14716 19312 14720
rect 19248 14660 19252 14716
rect 19252 14660 19308 14716
rect 19308 14660 19312 14716
rect 19248 14656 19312 14660
rect 19328 14716 19392 14720
rect 19328 14660 19332 14716
rect 19332 14660 19388 14716
rect 19388 14660 19392 14716
rect 19328 14656 19392 14660
rect 19408 14716 19472 14720
rect 19408 14660 19412 14716
rect 19412 14660 19468 14716
rect 19468 14660 19472 14716
rect 19408 14656 19472 14660
rect 5506 14172 5570 14176
rect 5506 14116 5510 14172
rect 5510 14116 5566 14172
rect 5566 14116 5570 14172
rect 5506 14112 5570 14116
rect 5586 14172 5650 14176
rect 5586 14116 5590 14172
rect 5590 14116 5646 14172
rect 5646 14116 5650 14172
rect 5586 14112 5650 14116
rect 5666 14172 5730 14176
rect 5666 14116 5670 14172
rect 5670 14116 5726 14172
rect 5726 14116 5730 14172
rect 5666 14112 5730 14116
rect 5746 14172 5810 14176
rect 5746 14116 5750 14172
rect 5750 14116 5806 14172
rect 5806 14116 5810 14172
rect 5746 14112 5810 14116
rect 14614 14172 14678 14176
rect 14614 14116 14618 14172
rect 14618 14116 14674 14172
rect 14674 14116 14678 14172
rect 14614 14112 14678 14116
rect 14694 14172 14758 14176
rect 14694 14116 14698 14172
rect 14698 14116 14754 14172
rect 14754 14116 14758 14172
rect 14694 14112 14758 14116
rect 14774 14172 14838 14176
rect 14774 14116 14778 14172
rect 14778 14116 14834 14172
rect 14834 14116 14838 14172
rect 14774 14112 14838 14116
rect 14854 14172 14918 14176
rect 14854 14116 14858 14172
rect 14858 14116 14914 14172
rect 14914 14116 14918 14172
rect 14854 14112 14918 14116
rect 23722 14172 23786 14176
rect 23722 14116 23726 14172
rect 23726 14116 23782 14172
rect 23782 14116 23786 14172
rect 23722 14112 23786 14116
rect 23802 14172 23866 14176
rect 23802 14116 23806 14172
rect 23806 14116 23862 14172
rect 23862 14116 23866 14172
rect 23802 14112 23866 14116
rect 23882 14172 23946 14176
rect 23882 14116 23886 14172
rect 23886 14116 23942 14172
rect 23942 14116 23946 14172
rect 23882 14112 23946 14116
rect 23962 14172 24026 14176
rect 23962 14116 23966 14172
rect 23966 14116 24022 14172
rect 24022 14116 24026 14172
rect 23962 14112 24026 14116
rect 10060 13628 10124 13632
rect 10060 13572 10064 13628
rect 10064 13572 10120 13628
rect 10120 13572 10124 13628
rect 10060 13568 10124 13572
rect 10140 13628 10204 13632
rect 10140 13572 10144 13628
rect 10144 13572 10200 13628
rect 10200 13572 10204 13628
rect 10140 13568 10204 13572
rect 10220 13628 10284 13632
rect 10220 13572 10224 13628
rect 10224 13572 10280 13628
rect 10280 13572 10284 13628
rect 10220 13568 10284 13572
rect 10300 13628 10364 13632
rect 10300 13572 10304 13628
rect 10304 13572 10360 13628
rect 10360 13572 10364 13628
rect 10300 13568 10364 13572
rect 19168 13628 19232 13632
rect 19168 13572 19172 13628
rect 19172 13572 19228 13628
rect 19228 13572 19232 13628
rect 19168 13568 19232 13572
rect 19248 13628 19312 13632
rect 19248 13572 19252 13628
rect 19252 13572 19308 13628
rect 19308 13572 19312 13628
rect 19248 13568 19312 13572
rect 19328 13628 19392 13632
rect 19328 13572 19332 13628
rect 19332 13572 19388 13628
rect 19388 13572 19392 13628
rect 19328 13568 19392 13572
rect 19408 13628 19472 13632
rect 19408 13572 19412 13628
rect 19412 13572 19468 13628
rect 19468 13572 19472 13628
rect 19408 13568 19472 13572
rect 5506 13084 5570 13088
rect 5506 13028 5510 13084
rect 5510 13028 5566 13084
rect 5566 13028 5570 13084
rect 5506 13024 5570 13028
rect 5586 13084 5650 13088
rect 5586 13028 5590 13084
rect 5590 13028 5646 13084
rect 5646 13028 5650 13084
rect 5586 13024 5650 13028
rect 5666 13084 5730 13088
rect 5666 13028 5670 13084
rect 5670 13028 5726 13084
rect 5726 13028 5730 13084
rect 5666 13024 5730 13028
rect 5746 13084 5810 13088
rect 5746 13028 5750 13084
rect 5750 13028 5806 13084
rect 5806 13028 5810 13084
rect 5746 13024 5810 13028
rect 14614 13084 14678 13088
rect 14614 13028 14618 13084
rect 14618 13028 14674 13084
rect 14674 13028 14678 13084
rect 14614 13024 14678 13028
rect 14694 13084 14758 13088
rect 14694 13028 14698 13084
rect 14698 13028 14754 13084
rect 14754 13028 14758 13084
rect 14694 13024 14758 13028
rect 14774 13084 14838 13088
rect 14774 13028 14778 13084
rect 14778 13028 14834 13084
rect 14834 13028 14838 13084
rect 14774 13024 14838 13028
rect 14854 13084 14918 13088
rect 14854 13028 14858 13084
rect 14858 13028 14914 13084
rect 14914 13028 14918 13084
rect 14854 13024 14918 13028
rect 23722 13084 23786 13088
rect 23722 13028 23726 13084
rect 23726 13028 23782 13084
rect 23782 13028 23786 13084
rect 23722 13024 23786 13028
rect 23802 13084 23866 13088
rect 23802 13028 23806 13084
rect 23806 13028 23862 13084
rect 23862 13028 23866 13084
rect 23802 13024 23866 13028
rect 23882 13084 23946 13088
rect 23882 13028 23886 13084
rect 23886 13028 23942 13084
rect 23942 13028 23946 13084
rect 23882 13024 23946 13028
rect 23962 13084 24026 13088
rect 23962 13028 23966 13084
rect 23966 13028 24022 13084
rect 24022 13028 24026 13084
rect 23962 13024 24026 13028
rect 10060 12540 10124 12544
rect 10060 12484 10064 12540
rect 10064 12484 10120 12540
rect 10120 12484 10124 12540
rect 10060 12480 10124 12484
rect 10140 12540 10204 12544
rect 10140 12484 10144 12540
rect 10144 12484 10200 12540
rect 10200 12484 10204 12540
rect 10140 12480 10204 12484
rect 10220 12540 10284 12544
rect 10220 12484 10224 12540
rect 10224 12484 10280 12540
rect 10280 12484 10284 12540
rect 10220 12480 10284 12484
rect 10300 12540 10364 12544
rect 10300 12484 10304 12540
rect 10304 12484 10360 12540
rect 10360 12484 10364 12540
rect 10300 12480 10364 12484
rect 19168 12540 19232 12544
rect 19168 12484 19172 12540
rect 19172 12484 19228 12540
rect 19228 12484 19232 12540
rect 19168 12480 19232 12484
rect 19248 12540 19312 12544
rect 19248 12484 19252 12540
rect 19252 12484 19308 12540
rect 19308 12484 19312 12540
rect 19248 12480 19312 12484
rect 19328 12540 19392 12544
rect 19328 12484 19332 12540
rect 19332 12484 19388 12540
rect 19388 12484 19392 12540
rect 19328 12480 19392 12484
rect 19408 12540 19472 12544
rect 19408 12484 19412 12540
rect 19412 12484 19468 12540
rect 19468 12484 19472 12540
rect 19408 12480 19472 12484
rect 5506 11996 5570 12000
rect 5506 11940 5510 11996
rect 5510 11940 5566 11996
rect 5566 11940 5570 11996
rect 5506 11936 5570 11940
rect 5586 11996 5650 12000
rect 5586 11940 5590 11996
rect 5590 11940 5646 11996
rect 5646 11940 5650 11996
rect 5586 11936 5650 11940
rect 5666 11996 5730 12000
rect 5666 11940 5670 11996
rect 5670 11940 5726 11996
rect 5726 11940 5730 11996
rect 5666 11936 5730 11940
rect 5746 11996 5810 12000
rect 5746 11940 5750 11996
rect 5750 11940 5806 11996
rect 5806 11940 5810 11996
rect 5746 11936 5810 11940
rect 14614 11996 14678 12000
rect 14614 11940 14618 11996
rect 14618 11940 14674 11996
rect 14674 11940 14678 11996
rect 14614 11936 14678 11940
rect 14694 11996 14758 12000
rect 14694 11940 14698 11996
rect 14698 11940 14754 11996
rect 14754 11940 14758 11996
rect 14694 11936 14758 11940
rect 14774 11996 14838 12000
rect 14774 11940 14778 11996
rect 14778 11940 14834 11996
rect 14834 11940 14838 11996
rect 14774 11936 14838 11940
rect 14854 11996 14918 12000
rect 14854 11940 14858 11996
rect 14858 11940 14914 11996
rect 14914 11940 14918 11996
rect 14854 11936 14918 11940
rect 23722 11996 23786 12000
rect 23722 11940 23726 11996
rect 23726 11940 23782 11996
rect 23782 11940 23786 11996
rect 23722 11936 23786 11940
rect 23802 11996 23866 12000
rect 23802 11940 23806 11996
rect 23806 11940 23862 11996
rect 23862 11940 23866 11996
rect 23802 11936 23866 11940
rect 23882 11996 23946 12000
rect 23882 11940 23886 11996
rect 23886 11940 23942 11996
rect 23942 11940 23946 11996
rect 23882 11936 23946 11940
rect 23962 11996 24026 12000
rect 23962 11940 23966 11996
rect 23966 11940 24022 11996
rect 24022 11940 24026 11996
rect 23962 11936 24026 11940
rect 10060 11452 10124 11456
rect 10060 11396 10064 11452
rect 10064 11396 10120 11452
rect 10120 11396 10124 11452
rect 10060 11392 10124 11396
rect 10140 11452 10204 11456
rect 10140 11396 10144 11452
rect 10144 11396 10200 11452
rect 10200 11396 10204 11452
rect 10140 11392 10204 11396
rect 10220 11452 10284 11456
rect 10220 11396 10224 11452
rect 10224 11396 10280 11452
rect 10280 11396 10284 11452
rect 10220 11392 10284 11396
rect 10300 11452 10364 11456
rect 10300 11396 10304 11452
rect 10304 11396 10360 11452
rect 10360 11396 10364 11452
rect 10300 11392 10364 11396
rect 19168 11452 19232 11456
rect 19168 11396 19172 11452
rect 19172 11396 19228 11452
rect 19228 11396 19232 11452
rect 19168 11392 19232 11396
rect 19248 11452 19312 11456
rect 19248 11396 19252 11452
rect 19252 11396 19308 11452
rect 19308 11396 19312 11452
rect 19248 11392 19312 11396
rect 19328 11452 19392 11456
rect 19328 11396 19332 11452
rect 19332 11396 19388 11452
rect 19388 11396 19392 11452
rect 19328 11392 19392 11396
rect 19408 11452 19472 11456
rect 19408 11396 19412 11452
rect 19412 11396 19468 11452
rect 19468 11396 19472 11452
rect 19408 11392 19472 11396
rect 10916 11052 10980 11116
rect 5506 10908 5570 10912
rect 5506 10852 5510 10908
rect 5510 10852 5566 10908
rect 5566 10852 5570 10908
rect 5506 10848 5570 10852
rect 5586 10908 5650 10912
rect 5586 10852 5590 10908
rect 5590 10852 5646 10908
rect 5646 10852 5650 10908
rect 5586 10848 5650 10852
rect 5666 10908 5730 10912
rect 5666 10852 5670 10908
rect 5670 10852 5726 10908
rect 5726 10852 5730 10908
rect 5666 10848 5730 10852
rect 5746 10908 5810 10912
rect 5746 10852 5750 10908
rect 5750 10852 5806 10908
rect 5806 10852 5810 10908
rect 5746 10848 5810 10852
rect 14614 10908 14678 10912
rect 14614 10852 14618 10908
rect 14618 10852 14674 10908
rect 14674 10852 14678 10908
rect 14614 10848 14678 10852
rect 14694 10908 14758 10912
rect 14694 10852 14698 10908
rect 14698 10852 14754 10908
rect 14754 10852 14758 10908
rect 14694 10848 14758 10852
rect 14774 10908 14838 10912
rect 14774 10852 14778 10908
rect 14778 10852 14834 10908
rect 14834 10852 14838 10908
rect 14774 10848 14838 10852
rect 14854 10908 14918 10912
rect 14854 10852 14858 10908
rect 14858 10852 14914 10908
rect 14914 10852 14918 10908
rect 14854 10848 14918 10852
rect 23722 10908 23786 10912
rect 23722 10852 23726 10908
rect 23726 10852 23782 10908
rect 23782 10852 23786 10908
rect 23722 10848 23786 10852
rect 23802 10908 23866 10912
rect 23802 10852 23806 10908
rect 23806 10852 23862 10908
rect 23862 10852 23866 10908
rect 23802 10848 23866 10852
rect 23882 10908 23946 10912
rect 23882 10852 23886 10908
rect 23886 10852 23942 10908
rect 23942 10852 23946 10908
rect 23882 10848 23946 10852
rect 23962 10908 24026 10912
rect 23962 10852 23966 10908
rect 23966 10852 24022 10908
rect 24022 10852 24026 10908
rect 23962 10848 24026 10852
rect 10060 10364 10124 10368
rect 10060 10308 10064 10364
rect 10064 10308 10120 10364
rect 10120 10308 10124 10364
rect 10060 10304 10124 10308
rect 10140 10364 10204 10368
rect 10140 10308 10144 10364
rect 10144 10308 10200 10364
rect 10200 10308 10204 10364
rect 10140 10304 10204 10308
rect 10220 10364 10284 10368
rect 10220 10308 10224 10364
rect 10224 10308 10280 10364
rect 10280 10308 10284 10364
rect 10220 10304 10284 10308
rect 10300 10364 10364 10368
rect 10300 10308 10304 10364
rect 10304 10308 10360 10364
rect 10360 10308 10364 10364
rect 10300 10304 10364 10308
rect 19168 10364 19232 10368
rect 19168 10308 19172 10364
rect 19172 10308 19228 10364
rect 19228 10308 19232 10364
rect 19168 10304 19232 10308
rect 19248 10364 19312 10368
rect 19248 10308 19252 10364
rect 19252 10308 19308 10364
rect 19308 10308 19312 10364
rect 19248 10304 19312 10308
rect 19328 10364 19392 10368
rect 19328 10308 19332 10364
rect 19332 10308 19388 10364
rect 19388 10308 19392 10364
rect 19328 10304 19392 10308
rect 19408 10364 19472 10368
rect 19408 10308 19412 10364
rect 19412 10308 19468 10364
rect 19468 10308 19472 10364
rect 19408 10304 19472 10308
rect 5506 9820 5570 9824
rect 5506 9764 5510 9820
rect 5510 9764 5566 9820
rect 5566 9764 5570 9820
rect 5506 9760 5570 9764
rect 5586 9820 5650 9824
rect 5586 9764 5590 9820
rect 5590 9764 5646 9820
rect 5646 9764 5650 9820
rect 5586 9760 5650 9764
rect 5666 9820 5730 9824
rect 5666 9764 5670 9820
rect 5670 9764 5726 9820
rect 5726 9764 5730 9820
rect 5666 9760 5730 9764
rect 5746 9820 5810 9824
rect 5746 9764 5750 9820
rect 5750 9764 5806 9820
rect 5806 9764 5810 9820
rect 5746 9760 5810 9764
rect 14614 9820 14678 9824
rect 14614 9764 14618 9820
rect 14618 9764 14674 9820
rect 14674 9764 14678 9820
rect 14614 9760 14678 9764
rect 14694 9820 14758 9824
rect 14694 9764 14698 9820
rect 14698 9764 14754 9820
rect 14754 9764 14758 9820
rect 14694 9760 14758 9764
rect 14774 9820 14838 9824
rect 14774 9764 14778 9820
rect 14778 9764 14834 9820
rect 14834 9764 14838 9820
rect 14774 9760 14838 9764
rect 14854 9820 14918 9824
rect 14854 9764 14858 9820
rect 14858 9764 14914 9820
rect 14914 9764 14918 9820
rect 14854 9760 14918 9764
rect 23722 9820 23786 9824
rect 23722 9764 23726 9820
rect 23726 9764 23782 9820
rect 23782 9764 23786 9820
rect 23722 9760 23786 9764
rect 23802 9820 23866 9824
rect 23802 9764 23806 9820
rect 23806 9764 23862 9820
rect 23862 9764 23866 9820
rect 23802 9760 23866 9764
rect 23882 9820 23946 9824
rect 23882 9764 23886 9820
rect 23886 9764 23942 9820
rect 23942 9764 23946 9820
rect 23882 9760 23946 9764
rect 23962 9820 24026 9824
rect 23962 9764 23966 9820
rect 23966 9764 24022 9820
rect 24022 9764 24026 9820
rect 23962 9760 24026 9764
rect 9812 9420 9876 9484
rect 10060 9276 10124 9280
rect 10060 9220 10064 9276
rect 10064 9220 10120 9276
rect 10120 9220 10124 9276
rect 10060 9216 10124 9220
rect 10140 9276 10204 9280
rect 10140 9220 10144 9276
rect 10144 9220 10200 9276
rect 10200 9220 10204 9276
rect 10140 9216 10204 9220
rect 10220 9276 10284 9280
rect 10220 9220 10224 9276
rect 10224 9220 10280 9276
rect 10280 9220 10284 9276
rect 10220 9216 10284 9220
rect 10300 9276 10364 9280
rect 10300 9220 10304 9276
rect 10304 9220 10360 9276
rect 10360 9220 10364 9276
rect 10300 9216 10364 9220
rect 19168 9276 19232 9280
rect 19168 9220 19172 9276
rect 19172 9220 19228 9276
rect 19228 9220 19232 9276
rect 19168 9216 19232 9220
rect 19248 9276 19312 9280
rect 19248 9220 19252 9276
rect 19252 9220 19308 9276
rect 19308 9220 19312 9276
rect 19248 9216 19312 9220
rect 19328 9276 19392 9280
rect 19328 9220 19332 9276
rect 19332 9220 19388 9276
rect 19388 9220 19392 9276
rect 19328 9216 19392 9220
rect 19408 9276 19472 9280
rect 19408 9220 19412 9276
rect 19412 9220 19468 9276
rect 19468 9220 19472 9276
rect 19408 9216 19472 9220
rect 5506 8732 5570 8736
rect 5506 8676 5510 8732
rect 5510 8676 5566 8732
rect 5566 8676 5570 8732
rect 5506 8672 5570 8676
rect 5586 8732 5650 8736
rect 5586 8676 5590 8732
rect 5590 8676 5646 8732
rect 5646 8676 5650 8732
rect 5586 8672 5650 8676
rect 5666 8732 5730 8736
rect 5666 8676 5670 8732
rect 5670 8676 5726 8732
rect 5726 8676 5730 8732
rect 5666 8672 5730 8676
rect 5746 8732 5810 8736
rect 5746 8676 5750 8732
rect 5750 8676 5806 8732
rect 5806 8676 5810 8732
rect 5746 8672 5810 8676
rect 14614 8732 14678 8736
rect 14614 8676 14618 8732
rect 14618 8676 14674 8732
rect 14674 8676 14678 8732
rect 14614 8672 14678 8676
rect 14694 8732 14758 8736
rect 14694 8676 14698 8732
rect 14698 8676 14754 8732
rect 14754 8676 14758 8732
rect 14694 8672 14758 8676
rect 14774 8732 14838 8736
rect 14774 8676 14778 8732
rect 14778 8676 14834 8732
rect 14834 8676 14838 8732
rect 14774 8672 14838 8676
rect 14854 8732 14918 8736
rect 14854 8676 14858 8732
rect 14858 8676 14914 8732
rect 14914 8676 14918 8732
rect 14854 8672 14918 8676
rect 23722 8732 23786 8736
rect 23722 8676 23726 8732
rect 23726 8676 23782 8732
rect 23782 8676 23786 8732
rect 23722 8672 23786 8676
rect 23802 8732 23866 8736
rect 23802 8676 23806 8732
rect 23806 8676 23862 8732
rect 23862 8676 23866 8732
rect 23802 8672 23866 8676
rect 23882 8732 23946 8736
rect 23882 8676 23886 8732
rect 23886 8676 23942 8732
rect 23942 8676 23946 8732
rect 23882 8672 23946 8676
rect 23962 8732 24026 8736
rect 23962 8676 23966 8732
rect 23966 8676 24022 8732
rect 24022 8676 24026 8732
rect 23962 8672 24026 8676
rect 10060 8188 10124 8192
rect 10060 8132 10064 8188
rect 10064 8132 10120 8188
rect 10120 8132 10124 8188
rect 10060 8128 10124 8132
rect 10140 8188 10204 8192
rect 10140 8132 10144 8188
rect 10144 8132 10200 8188
rect 10200 8132 10204 8188
rect 10140 8128 10204 8132
rect 10220 8188 10284 8192
rect 10220 8132 10224 8188
rect 10224 8132 10280 8188
rect 10280 8132 10284 8188
rect 10220 8128 10284 8132
rect 10300 8188 10364 8192
rect 10300 8132 10304 8188
rect 10304 8132 10360 8188
rect 10360 8132 10364 8188
rect 10300 8128 10364 8132
rect 19168 8188 19232 8192
rect 19168 8132 19172 8188
rect 19172 8132 19228 8188
rect 19228 8132 19232 8188
rect 19168 8128 19232 8132
rect 19248 8188 19312 8192
rect 19248 8132 19252 8188
rect 19252 8132 19308 8188
rect 19308 8132 19312 8188
rect 19248 8128 19312 8132
rect 19328 8188 19392 8192
rect 19328 8132 19332 8188
rect 19332 8132 19388 8188
rect 19388 8132 19392 8188
rect 19328 8128 19392 8132
rect 19408 8188 19472 8192
rect 19408 8132 19412 8188
rect 19412 8132 19468 8188
rect 19468 8132 19472 8188
rect 19408 8128 19472 8132
rect 5506 7644 5570 7648
rect 5506 7588 5510 7644
rect 5510 7588 5566 7644
rect 5566 7588 5570 7644
rect 5506 7584 5570 7588
rect 5586 7644 5650 7648
rect 5586 7588 5590 7644
rect 5590 7588 5646 7644
rect 5646 7588 5650 7644
rect 5586 7584 5650 7588
rect 5666 7644 5730 7648
rect 5666 7588 5670 7644
rect 5670 7588 5726 7644
rect 5726 7588 5730 7644
rect 5666 7584 5730 7588
rect 5746 7644 5810 7648
rect 5746 7588 5750 7644
rect 5750 7588 5806 7644
rect 5806 7588 5810 7644
rect 5746 7584 5810 7588
rect 14614 7644 14678 7648
rect 14614 7588 14618 7644
rect 14618 7588 14674 7644
rect 14674 7588 14678 7644
rect 14614 7584 14678 7588
rect 14694 7644 14758 7648
rect 14694 7588 14698 7644
rect 14698 7588 14754 7644
rect 14754 7588 14758 7644
rect 14694 7584 14758 7588
rect 14774 7644 14838 7648
rect 14774 7588 14778 7644
rect 14778 7588 14834 7644
rect 14834 7588 14838 7644
rect 14774 7584 14838 7588
rect 14854 7644 14918 7648
rect 14854 7588 14858 7644
rect 14858 7588 14914 7644
rect 14914 7588 14918 7644
rect 14854 7584 14918 7588
rect 23722 7644 23786 7648
rect 23722 7588 23726 7644
rect 23726 7588 23782 7644
rect 23782 7588 23786 7644
rect 23722 7584 23786 7588
rect 23802 7644 23866 7648
rect 23802 7588 23806 7644
rect 23806 7588 23862 7644
rect 23862 7588 23866 7644
rect 23802 7584 23866 7588
rect 23882 7644 23946 7648
rect 23882 7588 23886 7644
rect 23886 7588 23942 7644
rect 23942 7588 23946 7644
rect 23882 7584 23946 7588
rect 23962 7644 24026 7648
rect 23962 7588 23966 7644
rect 23966 7588 24022 7644
rect 24022 7588 24026 7644
rect 23962 7584 24026 7588
rect 10060 7100 10124 7104
rect 10060 7044 10064 7100
rect 10064 7044 10120 7100
rect 10120 7044 10124 7100
rect 10060 7040 10124 7044
rect 10140 7100 10204 7104
rect 10140 7044 10144 7100
rect 10144 7044 10200 7100
rect 10200 7044 10204 7100
rect 10140 7040 10204 7044
rect 10220 7100 10284 7104
rect 10220 7044 10224 7100
rect 10224 7044 10280 7100
rect 10280 7044 10284 7100
rect 10220 7040 10284 7044
rect 10300 7100 10364 7104
rect 10300 7044 10304 7100
rect 10304 7044 10360 7100
rect 10360 7044 10364 7100
rect 10300 7040 10364 7044
rect 19168 7100 19232 7104
rect 19168 7044 19172 7100
rect 19172 7044 19228 7100
rect 19228 7044 19232 7100
rect 19168 7040 19232 7044
rect 19248 7100 19312 7104
rect 19248 7044 19252 7100
rect 19252 7044 19308 7100
rect 19308 7044 19312 7100
rect 19248 7040 19312 7044
rect 19328 7100 19392 7104
rect 19328 7044 19332 7100
rect 19332 7044 19388 7100
rect 19388 7044 19392 7100
rect 19328 7040 19392 7044
rect 19408 7100 19472 7104
rect 19408 7044 19412 7100
rect 19412 7044 19468 7100
rect 19468 7044 19472 7100
rect 19408 7040 19472 7044
rect 5506 6556 5570 6560
rect 5506 6500 5510 6556
rect 5510 6500 5566 6556
rect 5566 6500 5570 6556
rect 5506 6496 5570 6500
rect 5586 6556 5650 6560
rect 5586 6500 5590 6556
rect 5590 6500 5646 6556
rect 5646 6500 5650 6556
rect 5586 6496 5650 6500
rect 5666 6556 5730 6560
rect 5666 6500 5670 6556
rect 5670 6500 5726 6556
rect 5726 6500 5730 6556
rect 5666 6496 5730 6500
rect 5746 6556 5810 6560
rect 5746 6500 5750 6556
rect 5750 6500 5806 6556
rect 5806 6500 5810 6556
rect 5746 6496 5810 6500
rect 14614 6556 14678 6560
rect 14614 6500 14618 6556
rect 14618 6500 14674 6556
rect 14674 6500 14678 6556
rect 14614 6496 14678 6500
rect 14694 6556 14758 6560
rect 14694 6500 14698 6556
rect 14698 6500 14754 6556
rect 14754 6500 14758 6556
rect 14694 6496 14758 6500
rect 14774 6556 14838 6560
rect 14774 6500 14778 6556
rect 14778 6500 14834 6556
rect 14834 6500 14838 6556
rect 14774 6496 14838 6500
rect 14854 6556 14918 6560
rect 14854 6500 14858 6556
rect 14858 6500 14914 6556
rect 14914 6500 14918 6556
rect 14854 6496 14918 6500
rect 23722 6556 23786 6560
rect 23722 6500 23726 6556
rect 23726 6500 23782 6556
rect 23782 6500 23786 6556
rect 23722 6496 23786 6500
rect 23802 6556 23866 6560
rect 23802 6500 23806 6556
rect 23806 6500 23862 6556
rect 23862 6500 23866 6556
rect 23802 6496 23866 6500
rect 23882 6556 23946 6560
rect 23882 6500 23886 6556
rect 23886 6500 23942 6556
rect 23942 6500 23946 6556
rect 23882 6496 23946 6500
rect 23962 6556 24026 6560
rect 23962 6500 23966 6556
rect 23966 6500 24022 6556
rect 24022 6500 24026 6556
rect 23962 6496 24026 6500
rect 10060 6012 10124 6016
rect 10060 5956 10064 6012
rect 10064 5956 10120 6012
rect 10120 5956 10124 6012
rect 10060 5952 10124 5956
rect 10140 6012 10204 6016
rect 10140 5956 10144 6012
rect 10144 5956 10200 6012
rect 10200 5956 10204 6012
rect 10140 5952 10204 5956
rect 10220 6012 10284 6016
rect 10220 5956 10224 6012
rect 10224 5956 10280 6012
rect 10280 5956 10284 6012
rect 10220 5952 10284 5956
rect 10300 6012 10364 6016
rect 10300 5956 10304 6012
rect 10304 5956 10360 6012
rect 10360 5956 10364 6012
rect 10300 5952 10364 5956
rect 19168 6012 19232 6016
rect 19168 5956 19172 6012
rect 19172 5956 19228 6012
rect 19228 5956 19232 6012
rect 19168 5952 19232 5956
rect 19248 6012 19312 6016
rect 19248 5956 19252 6012
rect 19252 5956 19308 6012
rect 19308 5956 19312 6012
rect 19248 5952 19312 5956
rect 19328 6012 19392 6016
rect 19328 5956 19332 6012
rect 19332 5956 19388 6012
rect 19388 5956 19392 6012
rect 19328 5952 19392 5956
rect 19408 6012 19472 6016
rect 19408 5956 19412 6012
rect 19412 5956 19468 6012
rect 19468 5956 19472 6012
rect 19408 5952 19472 5956
rect 5506 5468 5570 5472
rect 5506 5412 5510 5468
rect 5510 5412 5566 5468
rect 5566 5412 5570 5468
rect 5506 5408 5570 5412
rect 5586 5468 5650 5472
rect 5586 5412 5590 5468
rect 5590 5412 5646 5468
rect 5646 5412 5650 5468
rect 5586 5408 5650 5412
rect 5666 5468 5730 5472
rect 5666 5412 5670 5468
rect 5670 5412 5726 5468
rect 5726 5412 5730 5468
rect 5666 5408 5730 5412
rect 5746 5468 5810 5472
rect 5746 5412 5750 5468
rect 5750 5412 5806 5468
rect 5806 5412 5810 5468
rect 5746 5408 5810 5412
rect 14614 5468 14678 5472
rect 14614 5412 14618 5468
rect 14618 5412 14674 5468
rect 14674 5412 14678 5468
rect 14614 5408 14678 5412
rect 14694 5468 14758 5472
rect 14694 5412 14698 5468
rect 14698 5412 14754 5468
rect 14754 5412 14758 5468
rect 14694 5408 14758 5412
rect 14774 5468 14838 5472
rect 14774 5412 14778 5468
rect 14778 5412 14834 5468
rect 14834 5412 14838 5468
rect 14774 5408 14838 5412
rect 14854 5468 14918 5472
rect 14854 5412 14858 5468
rect 14858 5412 14914 5468
rect 14914 5412 14918 5468
rect 14854 5408 14918 5412
rect 23722 5468 23786 5472
rect 23722 5412 23726 5468
rect 23726 5412 23782 5468
rect 23782 5412 23786 5468
rect 23722 5408 23786 5412
rect 23802 5468 23866 5472
rect 23802 5412 23806 5468
rect 23806 5412 23862 5468
rect 23862 5412 23866 5468
rect 23802 5408 23866 5412
rect 23882 5468 23946 5472
rect 23882 5412 23886 5468
rect 23886 5412 23942 5468
rect 23942 5412 23946 5468
rect 23882 5408 23946 5412
rect 23962 5468 24026 5472
rect 23962 5412 23966 5468
rect 23966 5412 24022 5468
rect 24022 5412 24026 5468
rect 23962 5408 24026 5412
rect 10060 4924 10124 4928
rect 10060 4868 10064 4924
rect 10064 4868 10120 4924
rect 10120 4868 10124 4924
rect 10060 4864 10124 4868
rect 10140 4924 10204 4928
rect 10140 4868 10144 4924
rect 10144 4868 10200 4924
rect 10200 4868 10204 4924
rect 10140 4864 10204 4868
rect 10220 4924 10284 4928
rect 10220 4868 10224 4924
rect 10224 4868 10280 4924
rect 10280 4868 10284 4924
rect 10220 4864 10284 4868
rect 10300 4924 10364 4928
rect 10300 4868 10304 4924
rect 10304 4868 10360 4924
rect 10360 4868 10364 4924
rect 10300 4864 10364 4868
rect 19168 4924 19232 4928
rect 19168 4868 19172 4924
rect 19172 4868 19228 4924
rect 19228 4868 19232 4924
rect 19168 4864 19232 4868
rect 19248 4924 19312 4928
rect 19248 4868 19252 4924
rect 19252 4868 19308 4924
rect 19308 4868 19312 4924
rect 19248 4864 19312 4868
rect 19328 4924 19392 4928
rect 19328 4868 19332 4924
rect 19332 4868 19388 4924
rect 19388 4868 19392 4924
rect 19328 4864 19392 4868
rect 19408 4924 19472 4928
rect 19408 4868 19412 4924
rect 19412 4868 19468 4924
rect 19468 4868 19472 4924
rect 19408 4864 19472 4868
rect 5506 4380 5570 4384
rect 5506 4324 5510 4380
rect 5510 4324 5566 4380
rect 5566 4324 5570 4380
rect 5506 4320 5570 4324
rect 5586 4380 5650 4384
rect 5586 4324 5590 4380
rect 5590 4324 5646 4380
rect 5646 4324 5650 4380
rect 5586 4320 5650 4324
rect 5666 4380 5730 4384
rect 5666 4324 5670 4380
rect 5670 4324 5726 4380
rect 5726 4324 5730 4380
rect 5666 4320 5730 4324
rect 5746 4380 5810 4384
rect 5746 4324 5750 4380
rect 5750 4324 5806 4380
rect 5806 4324 5810 4380
rect 5746 4320 5810 4324
rect 14614 4380 14678 4384
rect 14614 4324 14618 4380
rect 14618 4324 14674 4380
rect 14674 4324 14678 4380
rect 14614 4320 14678 4324
rect 14694 4380 14758 4384
rect 14694 4324 14698 4380
rect 14698 4324 14754 4380
rect 14754 4324 14758 4380
rect 14694 4320 14758 4324
rect 14774 4380 14838 4384
rect 14774 4324 14778 4380
rect 14778 4324 14834 4380
rect 14834 4324 14838 4380
rect 14774 4320 14838 4324
rect 14854 4380 14918 4384
rect 14854 4324 14858 4380
rect 14858 4324 14914 4380
rect 14914 4324 14918 4380
rect 14854 4320 14918 4324
rect 23722 4380 23786 4384
rect 23722 4324 23726 4380
rect 23726 4324 23782 4380
rect 23782 4324 23786 4380
rect 23722 4320 23786 4324
rect 23802 4380 23866 4384
rect 23802 4324 23806 4380
rect 23806 4324 23862 4380
rect 23862 4324 23866 4380
rect 23802 4320 23866 4324
rect 23882 4380 23946 4384
rect 23882 4324 23886 4380
rect 23886 4324 23942 4380
rect 23942 4324 23946 4380
rect 23882 4320 23946 4324
rect 23962 4380 24026 4384
rect 23962 4324 23966 4380
rect 23966 4324 24022 4380
rect 24022 4324 24026 4380
rect 23962 4320 24026 4324
rect 26372 3980 26436 4044
rect 10060 3836 10124 3840
rect 10060 3780 10064 3836
rect 10064 3780 10120 3836
rect 10120 3780 10124 3836
rect 10060 3776 10124 3780
rect 10140 3836 10204 3840
rect 10140 3780 10144 3836
rect 10144 3780 10200 3836
rect 10200 3780 10204 3836
rect 10140 3776 10204 3780
rect 10220 3836 10284 3840
rect 10220 3780 10224 3836
rect 10224 3780 10280 3836
rect 10280 3780 10284 3836
rect 10220 3776 10284 3780
rect 10300 3836 10364 3840
rect 10300 3780 10304 3836
rect 10304 3780 10360 3836
rect 10360 3780 10364 3836
rect 10300 3776 10364 3780
rect 19168 3836 19232 3840
rect 19168 3780 19172 3836
rect 19172 3780 19228 3836
rect 19228 3780 19232 3836
rect 19168 3776 19232 3780
rect 19248 3836 19312 3840
rect 19248 3780 19252 3836
rect 19252 3780 19308 3836
rect 19308 3780 19312 3836
rect 19248 3776 19312 3780
rect 19328 3836 19392 3840
rect 19328 3780 19332 3836
rect 19332 3780 19388 3836
rect 19388 3780 19392 3836
rect 19328 3776 19392 3780
rect 19408 3836 19472 3840
rect 19408 3780 19412 3836
rect 19412 3780 19468 3836
rect 19468 3780 19472 3836
rect 19408 3776 19472 3780
rect 5506 3292 5570 3296
rect 5506 3236 5510 3292
rect 5510 3236 5566 3292
rect 5566 3236 5570 3292
rect 5506 3232 5570 3236
rect 5586 3292 5650 3296
rect 5586 3236 5590 3292
rect 5590 3236 5646 3292
rect 5646 3236 5650 3292
rect 5586 3232 5650 3236
rect 5666 3292 5730 3296
rect 5666 3236 5670 3292
rect 5670 3236 5726 3292
rect 5726 3236 5730 3292
rect 5666 3232 5730 3236
rect 5746 3292 5810 3296
rect 5746 3236 5750 3292
rect 5750 3236 5806 3292
rect 5806 3236 5810 3292
rect 5746 3232 5810 3236
rect 14614 3292 14678 3296
rect 14614 3236 14618 3292
rect 14618 3236 14674 3292
rect 14674 3236 14678 3292
rect 14614 3232 14678 3236
rect 14694 3292 14758 3296
rect 14694 3236 14698 3292
rect 14698 3236 14754 3292
rect 14754 3236 14758 3292
rect 14694 3232 14758 3236
rect 14774 3292 14838 3296
rect 14774 3236 14778 3292
rect 14778 3236 14834 3292
rect 14834 3236 14838 3292
rect 14774 3232 14838 3236
rect 14854 3292 14918 3296
rect 14854 3236 14858 3292
rect 14858 3236 14914 3292
rect 14914 3236 14918 3292
rect 14854 3232 14918 3236
rect 23722 3292 23786 3296
rect 23722 3236 23726 3292
rect 23726 3236 23782 3292
rect 23782 3236 23786 3292
rect 23722 3232 23786 3236
rect 23802 3292 23866 3296
rect 23802 3236 23806 3292
rect 23806 3236 23862 3292
rect 23862 3236 23866 3292
rect 23802 3232 23866 3236
rect 23882 3292 23946 3296
rect 23882 3236 23886 3292
rect 23886 3236 23942 3292
rect 23942 3236 23946 3292
rect 23882 3232 23946 3236
rect 23962 3292 24026 3296
rect 23962 3236 23966 3292
rect 23966 3236 24022 3292
rect 24022 3236 24026 3292
rect 23962 3232 24026 3236
rect 10060 2748 10124 2752
rect 10060 2692 10064 2748
rect 10064 2692 10120 2748
rect 10120 2692 10124 2748
rect 10060 2688 10124 2692
rect 10140 2748 10204 2752
rect 10140 2692 10144 2748
rect 10144 2692 10200 2748
rect 10200 2692 10204 2748
rect 10140 2688 10204 2692
rect 10220 2748 10284 2752
rect 10220 2692 10224 2748
rect 10224 2692 10280 2748
rect 10280 2692 10284 2748
rect 10220 2688 10284 2692
rect 10300 2748 10364 2752
rect 10300 2692 10304 2748
rect 10304 2692 10360 2748
rect 10360 2692 10364 2748
rect 10300 2688 10364 2692
rect 19168 2748 19232 2752
rect 19168 2692 19172 2748
rect 19172 2692 19228 2748
rect 19228 2692 19232 2748
rect 19168 2688 19232 2692
rect 19248 2748 19312 2752
rect 19248 2692 19252 2748
rect 19252 2692 19308 2748
rect 19308 2692 19312 2748
rect 19248 2688 19312 2692
rect 19328 2748 19392 2752
rect 19328 2692 19332 2748
rect 19332 2692 19388 2748
rect 19388 2692 19392 2748
rect 19328 2688 19392 2692
rect 19408 2748 19472 2752
rect 19408 2692 19412 2748
rect 19412 2692 19468 2748
rect 19468 2692 19472 2748
rect 19408 2688 19472 2692
rect 9812 2408 9876 2412
rect 9812 2352 9826 2408
rect 9826 2352 9876 2408
rect 9812 2348 9876 2352
rect 5506 2204 5570 2208
rect 5506 2148 5510 2204
rect 5510 2148 5566 2204
rect 5566 2148 5570 2204
rect 5506 2144 5570 2148
rect 5586 2204 5650 2208
rect 5586 2148 5590 2204
rect 5590 2148 5646 2204
rect 5646 2148 5650 2204
rect 5586 2144 5650 2148
rect 5666 2204 5730 2208
rect 5666 2148 5670 2204
rect 5670 2148 5726 2204
rect 5726 2148 5730 2204
rect 5666 2144 5730 2148
rect 5746 2204 5810 2208
rect 5746 2148 5750 2204
rect 5750 2148 5806 2204
rect 5806 2148 5810 2204
rect 5746 2144 5810 2148
rect 14614 2204 14678 2208
rect 14614 2148 14618 2204
rect 14618 2148 14674 2204
rect 14674 2148 14678 2204
rect 14614 2144 14678 2148
rect 14694 2204 14758 2208
rect 14694 2148 14698 2204
rect 14698 2148 14754 2204
rect 14754 2148 14758 2204
rect 14694 2144 14758 2148
rect 14774 2204 14838 2208
rect 14774 2148 14778 2204
rect 14778 2148 14834 2204
rect 14834 2148 14838 2204
rect 14774 2144 14838 2148
rect 14854 2204 14918 2208
rect 14854 2148 14858 2204
rect 14858 2148 14914 2204
rect 14914 2148 14918 2204
rect 14854 2144 14918 2148
rect 23722 2204 23786 2208
rect 23722 2148 23726 2204
rect 23726 2148 23782 2204
rect 23782 2148 23786 2204
rect 23722 2144 23786 2148
rect 23802 2204 23866 2208
rect 23802 2148 23806 2204
rect 23806 2148 23862 2204
rect 23862 2148 23866 2204
rect 23802 2144 23866 2148
rect 23882 2204 23946 2208
rect 23882 2148 23886 2204
rect 23886 2148 23942 2204
rect 23942 2148 23946 2204
rect 23882 2144 23946 2148
rect 23962 2204 24026 2208
rect 23962 2148 23966 2204
rect 23966 2148 24022 2204
rect 24022 2148 24026 2204
rect 23962 2144 24026 2148
<< metal4 >>
rect 5498 29408 5818 29424
rect 5498 29344 5506 29408
rect 5570 29344 5586 29408
rect 5650 29344 5666 29408
rect 5730 29344 5746 29408
rect 5810 29344 5818 29408
rect 5498 28320 5818 29344
rect 10052 28864 10372 29424
rect 10052 28800 10060 28864
rect 10124 28800 10140 28864
rect 10204 28800 10220 28864
rect 10284 28800 10300 28864
rect 10364 28800 10372 28864
rect 9811 28660 9877 28661
rect 9811 28596 9812 28660
rect 9876 28596 9877 28660
rect 9811 28595 9877 28596
rect 5498 28256 5506 28320
rect 5570 28256 5586 28320
rect 5650 28256 5666 28320
rect 5730 28256 5746 28320
rect 5810 28256 5818 28320
rect 5498 27232 5818 28256
rect 5498 27168 5506 27232
rect 5570 27168 5586 27232
rect 5650 27168 5666 27232
rect 5730 27168 5746 27232
rect 5810 27168 5818 27232
rect 5498 26144 5818 27168
rect 5498 26080 5506 26144
rect 5570 26080 5586 26144
rect 5650 26080 5666 26144
rect 5730 26080 5746 26144
rect 5810 26080 5818 26144
rect 5498 25056 5818 26080
rect 5498 24992 5506 25056
rect 5570 24992 5586 25056
rect 5650 24992 5666 25056
rect 5730 24992 5746 25056
rect 5810 24992 5818 25056
rect 5498 24912 5818 24992
rect 5498 24676 5540 24912
rect 5776 24676 5818 24912
rect 5498 23968 5818 24676
rect 9814 24173 9874 28595
rect 10052 27776 10372 28800
rect 10052 27712 10060 27776
rect 10124 27712 10140 27776
rect 10204 27712 10220 27776
rect 10284 27712 10300 27776
rect 10364 27712 10372 27776
rect 10052 26688 10372 27712
rect 10052 26624 10060 26688
rect 10124 26624 10140 26688
rect 10204 26624 10220 26688
rect 10284 26624 10300 26688
rect 10364 26624 10372 26688
rect 10052 25600 10372 26624
rect 10052 25536 10060 25600
rect 10124 25536 10140 25600
rect 10204 25536 10220 25600
rect 10284 25536 10300 25600
rect 10364 25536 10372 25600
rect 10052 24512 10372 25536
rect 10052 24448 10060 24512
rect 10124 24448 10140 24512
rect 10204 24448 10220 24512
rect 10284 24448 10300 24512
rect 10364 24448 10372 24512
rect 9811 24172 9877 24173
rect 9811 24108 9812 24172
rect 9876 24108 9877 24172
rect 9811 24107 9877 24108
rect 5498 23904 5506 23968
rect 5570 23904 5586 23968
rect 5650 23904 5666 23968
rect 5730 23904 5746 23968
rect 5810 23904 5818 23968
rect 5498 22880 5818 23904
rect 5498 22816 5506 22880
rect 5570 22816 5586 22880
rect 5650 22816 5666 22880
rect 5730 22816 5746 22880
rect 5810 22816 5818 22880
rect 5498 21792 5818 22816
rect 5498 21728 5506 21792
rect 5570 21728 5586 21792
rect 5650 21728 5666 21792
rect 5730 21728 5746 21792
rect 5810 21728 5818 21792
rect 5498 20704 5818 21728
rect 5498 20640 5506 20704
rect 5570 20640 5586 20704
rect 5650 20640 5666 20704
rect 5730 20640 5746 20704
rect 5810 20640 5818 20704
rect 5498 19616 5818 20640
rect 5498 19552 5506 19616
rect 5570 19552 5586 19616
rect 5650 19552 5666 19616
rect 5730 19552 5746 19616
rect 5810 19552 5818 19616
rect 5498 18528 5818 19552
rect 10052 23424 10372 24448
rect 10052 23360 10060 23424
rect 10124 23360 10140 23424
rect 10204 23360 10220 23424
rect 10284 23360 10300 23424
rect 10364 23360 10372 23424
rect 10052 22336 10372 23360
rect 10052 22272 10060 22336
rect 10124 22272 10140 22336
rect 10204 22272 10220 22336
rect 10284 22272 10300 22336
rect 10364 22272 10372 22336
rect 10052 21248 10372 22272
rect 10052 21184 10060 21248
rect 10124 21184 10140 21248
rect 10204 21184 10220 21248
rect 10284 21184 10300 21248
rect 10364 21184 10372 21248
rect 10052 20379 10372 21184
rect 10052 20160 10094 20379
rect 10330 20160 10372 20379
rect 10052 20096 10060 20160
rect 10124 20096 10140 20143
rect 10204 20096 10220 20143
rect 10284 20096 10300 20143
rect 10364 20096 10372 20160
rect 9811 19276 9877 19277
rect 9811 19212 9812 19276
rect 9876 19212 9877 19276
rect 9811 19211 9877 19212
rect 5498 18464 5506 18528
rect 5570 18464 5586 18528
rect 5650 18464 5666 18528
rect 5730 18464 5746 18528
rect 5810 18464 5818 18528
rect 5498 17440 5818 18464
rect 5498 17376 5506 17440
rect 5570 17376 5586 17440
rect 5650 17376 5666 17440
rect 5730 17376 5746 17440
rect 5810 17376 5818 17440
rect 5498 16352 5818 17376
rect 9814 17373 9874 19211
rect 10052 19072 10372 20096
rect 10052 19008 10060 19072
rect 10124 19008 10140 19072
rect 10204 19008 10220 19072
rect 10284 19008 10300 19072
rect 10364 19008 10372 19072
rect 10052 17984 10372 19008
rect 10052 17920 10060 17984
rect 10124 17920 10140 17984
rect 10204 17920 10220 17984
rect 10284 17920 10300 17984
rect 10364 17920 10372 17984
rect 9811 17372 9877 17373
rect 9811 17308 9812 17372
rect 9876 17308 9877 17372
rect 9811 17307 9877 17308
rect 5498 16288 5506 16352
rect 5570 16288 5586 16352
rect 5650 16288 5666 16352
rect 5730 16288 5746 16352
rect 5810 16288 5818 16352
rect 5498 15846 5818 16288
rect 5498 15610 5540 15846
rect 5776 15610 5818 15846
rect 5498 15264 5818 15610
rect 5498 15200 5506 15264
rect 5570 15200 5586 15264
rect 5650 15200 5666 15264
rect 5730 15200 5746 15264
rect 5810 15200 5818 15264
rect 5498 14176 5818 15200
rect 5498 14112 5506 14176
rect 5570 14112 5586 14176
rect 5650 14112 5666 14176
rect 5730 14112 5746 14176
rect 5810 14112 5818 14176
rect 5498 13088 5818 14112
rect 5498 13024 5506 13088
rect 5570 13024 5586 13088
rect 5650 13024 5666 13088
rect 5730 13024 5746 13088
rect 5810 13024 5818 13088
rect 5498 12000 5818 13024
rect 5498 11936 5506 12000
rect 5570 11936 5586 12000
rect 5650 11936 5666 12000
rect 5730 11936 5746 12000
rect 5810 11936 5818 12000
rect 5498 10912 5818 11936
rect 5498 10848 5506 10912
rect 5570 10848 5586 10912
rect 5650 10848 5666 10912
rect 5730 10848 5746 10912
rect 5810 10848 5818 10912
rect 5498 9824 5818 10848
rect 5498 9760 5506 9824
rect 5570 9760 5586 9824
rect 5650 9760 5666 9824
rect 5730 9760 5746 9824
rect 5810 9760 5818 9824
rect 5498 8736 5818 9760
rect 10052 16896 10372 17920
rect 10052 16832 10060 16896
rect 10124 16832 10140 16896
rect 10204 16832 10220 16896
rect 10284 16832 10300 16896
rect 10364 16832 10372 16896
rect 10052 15808 10372 16832
rect 14606 29408 14926 29424
rect 14606 29344 14614 29408
rect 14678 29344 14694 29408
rect 14758 29344 14774 29408
rect 14838 29344 14854 29408
rect 14918 29344 14926 29408
rect 14606 28320 14926 29344
rect 14606 28256 14614 28320
rect 14678 28256 14694 28320
rect 14758 28256 14774 28320
rect 14838 28256 14854 28320
rect 14918 28256 14926 28320
rect 14606 27232 14926 28256
rect 14606 27168 14614 27232
rect 14678 27168 14694 27232
rect 14758 27168 14774 27232
rect 14838 27168 14854 27232
rect 14918 27168 14926 27232
rect 14606 26144 14926 27168
rect 14606 26080 14614 26144
rect 14678 26080 14694 26144
rect 14758 26080 14774 26144
rect 14838 26080 14854 26144
rect 14918 26080 14926 26144
rect 14606 25056 14926 26080
rect 14606 24992 14614 25056
rect 14678 24992 14694 25056
rect 14758 24992 14774 25056
rect 14838 24992 14854 25056
rect 14918 24992 14926 25056
rect 14606 24912 14926 24992
rect 14606 24676 14648 24912
rect 14884 24676 14926 24912
rect 14606 23968 14926 24676
rect 14606 23904 14614 23968
rect 14678 23904 14694 23968
rect 14758 23904 14774 23968
rect 14838 23904 14854 23968
rect 14918 23904 14926 23968
rect 14606 22880 14926 23904
rect 14606 22816 14614 22880
rect 14678 22816 14694 22880
rect 14758 22816 14774 22880
rect 14838 22816 14854 22880
rect 14918 22816 14926 22880
rect 14606 21792 14926 22816
rect 14606 21728 14614 21792
rect 14678 21728 14694 21792
rect 14758 21728 14774 21792
rect 14838 21728 14854 21792
rect 14918 21728 14926 21792
rect 14606 20704 14926 21728
rect 14606 20640 14614 20704
rect 14678 20640 14694 20704
rect 14758 20640 14774 20704
rect 14838 20640 14854 20704
rect 14918 20640 14926 20704
rect 14606 19616 14926 20640
rect 14606 19552 14614 19616
rect 14678 19552 14694 19616
rect 14758 19552 14774 19616
rect 14838 19552 14854 19616
rect 14918 19552 14926 19616
rect 14606 18528 14926 19552
rect 14606 18464 14614 18528
rect 14678 18464 14694 18528
rect 14758 18464 14774 18528
rect 14838 18464 14854 18528
rect 14918 18464 14926 18528
rect 14606 17440 14926 18464
rect 14606 17376 14614 17440
rect 14678 17376 14694 17440
rect 14758 17376 14774 17440
rect 14838 17376 14854 17440
rect 14918 17376 14926 17440
rect 14606 16352 14926 17376
rect 14606 16288 14614 16352
rect 14678 16288 14694 16352
rect 14758 16288 14774 16352
rect 14838 16288 14854 16352
rect 14918 16288 14926 16352
rect 10915 16148 10981 16149
rect 10915 16084 10916 16148
rect 10980 16084 10981 16148
rect 10915 16083 10981 16084
rect 10052 15744 10060 15808
rect 10124 15744 10140 15808
rect 10204 15744 10220 15808
rect 10284 15744 10300 15808
rect 10364 15744 10372 15808
rect 10052 14720 10372 15744
rect 10052 14656 10060 14720
rect 10124 14656 10140 14720
rect 10204 14656 10220 14720
rect 10284 14656 10300 14720
rect 10364 14656 10372 14720
rect 10052 13632 10372 14656
rect 10052 13568 10060 13632
rect 10124 13568 10140 13632
rect 10204 13568 10220 13632
rect 10284 13568 10300 13632
rect 10364 13568 10372 13632
rect 10052 12544 10372 13568
rect 10052 12480 10060 12544
rect 10124 12480 10140 12544
rect 10204 12480 10220 12544
rect 10284 12480 10300 12544
rect 10364 12480 10372 12544
rect 10052 11456 10372 12480
rect 10052 11392 10060 11456
rect 10124 11392 10140 11456
rect 10204 11392 10220 11456
rect 10284 11392 10300 11456
rect 10364 11392 10372 11456
rect 10052 11312 10372 11392
rect 10052 11076 10094 11312
rect 10330 11076 10372 11312
rect 10918 11117 10978 16083
rect 14606 15846 14926 16288
rect 14606 15610 14648 15846
rect 14884 15610 14926 15846
rect 14606 15264 14926 15610
rect 14606 15200 14614 15264
rect 14678 15200 14694 15264
rect 14758 15200 14774 15264
rect 14838 15200 14854 15264
rect 14918 15200 14926 15264
rect 14606 14176 14926 15200
rect 14606 14112 14614 14176
rect 14678 14112 14694 14176
rect 14758 14112 14774 14176
rect 14838 14112 14854 14176
rect 14918 14112 14926 14176
rect 14606 13088 14926 14112
rect 14606 13024 14614 13088
rect 14678 13024 14694 13088
rect 14758 13024 14774 13088
rect 14838 13024 14854 13088
rect 14918 13024 14926 13088
rect 14606 12000 14926 13024
rect 14606 11936 14614 12000
rect 14678 11936 14694 12000
rect 14758 11936 14774 12000
rect 14838 11936 14854 12000
rect 14918 11936 14926 12000
rect 10052 10368 10372 11076
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 10052 10304 10060 10368
rect 10124 10304 10140 10368
rect 10204 10304 10220 10368
rect 10284 10304 10300 10368
rect 10364 10304 10372 10368
rect 9811 9484 9877 9485
rect 9811 9420 9812 9484
rect 9876 9420 9877 9484
rect 9811 9419 9877 9420
rect 5498 8672 5506 8736
rect 5570 8672 5586 8736
rect 5650 8672 5666 8736
rect 5730 8672 5746 8736
rect 5810 8672 5818 8736
rect 5498 7648 5818 8672
rect 5498 7584 5506 7648
rect 5570 7584 5586 7648
rect 5650 7584 5666 7648
rect 5730 7584 5746 7648
rect 5810 7584 5818 7648
rect 5498 6779 5818 7584
rect 5498 6560 5540 6779
rect 5776 6560 5818 6779
rect 5498 6496 5506 6560
rect 5570 6496 5586 6543
rect 5650 6496 5666 6543
rect 5730 6496 5746 6543
rect 5810 6496 5818 6560
rect 5498 5472 5818 6496
rect 5498 5408 5506 5472
rect 5570 5408 5586 5472
rect 5650 5408 5666 5472
rect 5730 5408 5746 5472
rect 5810 5408 5818 5472
rect 5498 4384 5818 5408
rect 5498 4320 5506 4384
rect 5570 4320 5586 4384
rect 5650 4320 5666 4384
rect 5730 4320 5746 4384
rect 5810 4320 5818 4384
rect 5498 3296 5818 4320
rect 5498 3232 5506 3296
rect 5570 3232 5586 3296
rect 5650 3232 5666 3296
rect 5730 3232 5746 3296
rect 5810 3232 5818 3296
rect 5498 2208 5818 3232
rect 9814 2413 9874 9419
rect 10052 9280 10372 10304
rect 10052 9216 10060 9280
rect 10124 9216 10140 9280
rect 10204 9216 10220 9280
rect 10284 9216 10300 9280
rect 10364 9216 10372 9280
rect 10052 8192 10372 9216
rect 10052 8128 10060 8192
rect 10124 8128 10140 8192
rect 10204 8128 10220 8192
rect 10284 8128 10300 8192
rect 10364 8128 10372 8192
rect 10052 7104 10372 8128
rect 10052 7040 10060 7104
rect 10124 7040 10140 7104
rect 10204 7040 10220 7104
rect 10284 7040 10300 7104
rect 10364 7040 10372 7104
rect 10052 6016 10372 7040
rect 10052 5952 10060 6016
rect 10124 5952 10140 6016
rect 10204 5952 10220 6016
rect 10284 5952 10300 6016
rect 10364 5952 10372 6016
rect 10052 4928 10372 5952
rect 10052 4864 10060 4928
rect 10124 4864 10140 4928
rect 10204 4864 10220 4928
rect 10284 4864 10300 4928
rect 10364 4864 10372 4928
rect 10052 3840 10372 4864
rect 10052 3776 10060 3840
rect 10124 3776 10140 3840
rect 10204 3776 10220 3840
rect 10284 3776 10300 3840
rect 10364 3776 10372 3840
rect 10052 2752 10372 3776
rect 10052 2688 10060 2752
rect 10124 2688 10140 2752
rect 10204 2688 10220 2752
rect 10284 2688 10300 2752
rect 10364 2688 10372 2752
rect 9811 2412 9877 2413
rect 9811 2348 9812 2412
rect 9876 2348 9877 2412
rect 9811 2347 9877 2348
rect 5498 2144 5506 2208
rect 5570 2144 5586 2208
rect 5650 2144 5666 2208
rect 5730 2144 5746 2208
rect 5810 2144 5818 2208
rect 5498 2128 5818 2144
rect 10052 2128 10372 2688
rect 14606 10912 14926 11936
rect 14606 10848 14614 10912
rect 14678 10848 14694 10912
rect 14758 10848 14774 10912
rect 14838 10848 14854 10912
rect 14918 10848 14926 10912
rect 14606 9824 14926 10848
rect 14606 9760 14614 9824
rect 14678 9760 14694 9824
rect 14758 9760 14774 9824
rect 14838 9760 14854 9824
rect 14918 9760 14926 9824
rect 14606 8736 14926 9760
rect 14606 8672 14614 8736
rect 14678 8672 14694 8736
rect 14758 8672 14774 8736
rect 14838 8672 14854 8736
rect 14918 8672 14926 8736
rect 14606 7648 14926 8672
rect 14606 7584 14614 7648
rect 14678 7584 14694 7648
rect 14758 7584 14774 7648
rect 14838 7584 14854 7648
rect 14918 7584 14926 7648
rect 14606 6779 14926 7584
rect 14606 6560 14648 6779
rect 14884 6560 14926 6779
rect 14606 6496 14614 6560
rect 14678 6496 14694 6543
rect 14758 6496 14774 6543
rect 14838 6496 14854 6543
rect 14918 6496 14926 6560
rect 14606 5472 14926 6496
rect 14606 5408 14614 5472
rect 14678 5408 14694 5472
rect 14758 5408 14774 5472
rect 14838 5408 14854 5472
rect 14918 5408 14926 5472
rect 14606 4384 14926 5408
rect 14606 4320 14614 4384
rect 14678 4320 14694 4384
rect 14758 4320 14774 4384
rect 14838 4320 14854 4384
rect 14918 4320 14926 4384
rect 14606 3296 14926 4320
rect 14606 3232 14614 3296
rect 14678 3232 14694 3296
rect 14758 3232 14774 3296
rect 14838 3232 14854 3296
rect 14918 3232 14926 3296
rect 14606 2208 14926 3232
rect 14606 2144 14614 2208
rect 14678 2144 14694 2208
rect 14758 2144 14774 2208
rect 14838 2144 14854 2208
rect 14918 2144 14926 2208
rect 14606 2128 14926 2144
rect 19160 28864 19480 29424
rect 19160 28800 19168 28864
rect 19232 28800 19248 28864
rect 19312 28800 19328 28864
rect 19392 28800 19408 28864
rect 19472 28800 19480 28864
rect 19160 27776 19480 28800
rect 19160 27712 19168 27776
rect 19232 27712 19248 27776
rect 19312 27712 19328 27776
rect 19392 27712 19408 27776
rect 19472 27712 19480 27776
rect 19160 26688 19480 27712
rect 19160 26624 19168 26688
rect 19232 26624 19248 26688
rect 19312 26624 19328 26688
rect 19392 26624 19408 26688
rect 19472 26624 19480 26688
rect 19160 25600 19480 26624
rect 19160 25536 19168 25600
rect 19232 25536 19248 25600
rect 19312 25536 19328 25600
rect 19392 25536 19408 25600
rect 19472 25536 19480 25600
rect 19160 24512 19480 25536
rect 19160 24448 19168 24512
rect 19232 24448 19248 24512
rect 19312 24448 19328 24512
rect 19392 24448 19408 24512
rect 19472 24448 19480 24512
rect 19160 23424 19480 24448
rect 19160 23360 19168 23424
rect 19232 23360 19248 23424
rect 19312 23360 19328 23424
rect 19392 23360 19408 23424
rect 19472 23360 19480 23424
rect 19160 22336 19480 23360
rect 19160 22272 19168 22336
rect 19232 22272 19248 22336
rect 19312 22272 19328 22336
rect 19392 22272 19408 22336
rect 19472 22272 19480 22336
rect 19160 21248 19480 22272
rect 19160 21184 19168 21248
rect 19232 21184 19248 21248
rect 19312 21184 19328 21248
rect 19392 21184 19408 21248
rect 19472 21184 19480 21248
rect 19160 20379 19480 21184
rect 19160 20160 19202 20379
rect 19438 20160 19480 20379
rect 19160 20096 19168 20160
rect 19232 20096 19248 20143
rect 19312 20096 19328 20143
rect 19392 20096 19408 20143
rect 19472 20096 19480 20160
rect 19160 19072 19480 20096
rect 19160 19008 19168 19072
rect 19232 19008 19248 19072
rect 19312 19008 19328 19072
rect 19392 19008 19408 19072
rect 19472 19008 19480 19072
rect 19160 17984 19480 19008
rect 19160 17920 19168 17984
rect 19232 17920 19248 17984
rect 19312 17920 19328 17984
rect 19392 17920 19408 17984
rect 19472 17920 19480 17984
rect 19160 16896 19480 17920
rect 19160 16832 19168 16896
rect 19232 16832 19248 16896
rect 19312 16832 19328 16896
rect 19392 16832 19408 16896
rect 19472 16832 19480 16896
rect 19160 15808 19480 16832
rect 19160 15744 19168 15808
rect 19232 15744 19248 15808
rect 19312 15744 19328 15808
rect 19392 15744 19408 15808
rect 19472 15744 19480 15808
rect 19160 14720 19480 15744
rect 19160 14656 19168 14720
rect 19232 14656 19248 14720
rect 19312 14656 19328 14720
rect 19392 14656 19408 14720
rect 19472 14656 19480 14720
rect 19160 13632 19480 14656
rect 19160 13568 19168 13632
rect 19232 13568 19248 13632
rect 19312 13568 19328 13632
rect 19392 13568 19408 13632
rect 19472 13568 19480 13632
rect 19160 12544 19480 13568
rect 19160 12480 19168 12544
rect 19232 12480 19248 12544
rect 19312 12480 19328 12544
rect 19392 12480 19408 12544
rect 19472 12480 19480 12544
rect 19160 11456 19480 12480
rect 19160 11392 19168 11456
rect 19232 11392 19248 11456
rect 19312 11392 19328 11456
rect 19392 11392 19408 11456
rect 19472 11392 19480 11456
rect 19160 11312 19480 11392
rect 19160 11076 19202 11312
rect 19438 11076 19480 11312
rect 19160 10368 19480 11076
rect 19160 10304 19168 10368
rect 19232 10304 19248 10368
rect 19312 10304 19328 10368
rect 19392 10304 19408 10368
rect 19472 10304 19480 10368
rect 19160 9280 19480 10304
rect 19160 9216 19168 9280
rect 19232 9216 19248 9280
rect 19312 9216 19328 9280
rect 19392 9216 19408 9280
rect 19472 9216 19480 9280
rect 19160 8192 19480 9216
rect 19160 8128 19168 8192
rect 19232 8128 19248 8192
rect 19312 8128 19328 8192
rect 19392 8128 19408 8192
rect 19472 8128 19480 8192
rect 19160 7104 19480 8128
rect 19160 7040 19168 7104
rect 19232 7040 19248 7104
rect 19312 7040 19328 7104
rect 19392 7040 19408 7104
rect 19472 7040 19480 7104
rect 19160 6016 19480 7040
rect 19160 5952 19168 6016
rect 19232 5952 19248 6016
rect 19312 5952 19328 6016
rect 19392 5952 19408 6016
rect 19472 5952 19480 6016
rect 19160 4928 19480 5952
rect 19160 4864 19168 4928
rect 19232 4864 19248 4928
rect 19312 4864 19328 4928
rect 19392 4864 19408 4928
rect 19472 4864 19480 4928
rect 19160 3840 19480 4864
rect 19160 3776 19168 3840
rect 19232 3776 19248 3840
rect 19312 3776 19328 3840
rect 19392 3776 19408 3840
rect 19472 3776 19480 3840
rect 19160 2752 19480 3776
rect 19160 2688 19168 2752
rect 19232 2688 19248 2752
rect 19312 2688 19328 2752
rect 19392 2688 19408 2752
rect 19472 2688 19480 2752
rect 19160 2128 19480 2688
rect 23714 29408 24034 29424
rect 23714 29344 23722 29408
rect 23786 29344 23802 29408
rect 23866 29344 23882 29408
rect 23946 29344 23962 29408
rect 24026 29344 24034 29408
rect 23714 28320 24034 29344
rect 23714 28256 23722 28320
rect 23786 28256 23802 28320
rect 23866 28256 23882 28320
rect 23946 28256 23962 28320
rect 24026 28256 24034 28320
rect 23714 27232 24034 28256
rect 23714 27168 23722 27232
rect 23786 27168 23802 27232
rect 23866 27168 23882 27232
rect 23946 27168 23962 27232
rect 24026 27168 24034 27232
rect 23714 26144 24034 27168
rect 23714 26080 23722 26144
rect 23786 26080 23802 26144
rect 23866 26080 23882 26144
rect 23946 26080 23962 26144
rect 24026 26080 24034 26144
rect 23714 25056 24034 26080
rect 23714 24992 23722 25056
rect 23786 24992 23802 25056
rect 23866 24992 23882 25056
rect 23946 24992 23962 25056
rect 24026 24992 24034 25056
rect 23714 24912 24034 24992
rect 23714 24676 23756 24912
rect 23992 24676 24034 24912
rect 23714 23968 24034 24676
rect 23714 23904 23722 23968
rect 23786 23904 23802 23968
rect 23866 23904 23882 23968
rect 23946 23904 23962 23968
rect 24026 23904 24034 23968
rect 23714 22880 24034 23904
rect 26371 23492 26437 23493
rect 26371 23428 26372 23492
rect 26436 23428 26437 23492
rect 26371 23427 26437 23428
rect 23714 22816 23722 22880
rect 23786 22816 23802 22880
rect 23866 22816 23882 22880
rect 23946 22816 23962 22880
rect 24026 22816 24034 22880
rect 23714 21792 24034 22816
rect 23714 21728 23722 21792
rect 23786 21728 23802 21792
rect 23866 21728 23882 21792
rect 23946 21728 23962 21792
rect 24026 21728 24034 21792
rect 23714 20704 24034 21728
rect 23714 20640 23722 20704
rect 23786 20640 23802 20704
rect 23866 20640 23882 20704
rect 23946 20640 23962 20704
rect 24026 20640 24034 20704
rect 23714 19616 24034 20640
rect 23714 19552 23722 19616
rect 23786 19552 23802 19616
rect 23866 19552 23882 19616
rect 23946 19552 23962 19616
rect 24026 19552 24034 19616
rect 23714 18528 24034 19552
rect 23714 18464 23722 18528
rect 23786 18464 23802 18528
rect 23866 18464 23882 18528
rect 23946 18464 23962 18528
rect 24026 18464 24034 18528
rect 23714 17440 24034 18464
rect 23714 17376 23722 17440
rect 23786 17376 23802 17440
rect 23866 17376 23882 17440
rect 23946 17376 23962 17440
rect 24026 17376 24034 17440
rect 23714 16352 24034 17376
rect 23714 16288 23722 16352
rect 23786 16288 23802 16352
rect 23866 16288 23882 16352
rect 23946 16288 23962 16352
rect 24026 16288 24034 16352
rect 23714 15846 24034 16288
rect 23714 15610 23756 15846
rect 23992 15610 24034 15846
rect 23714 15264 24034 15610
rect 23714 15200 23722 15264
rect 23786 15200 23802 15264
rect 23866 15200 23882 15264
rect 23946 15200 23962 15264
rect 24026 15200 24034 15264
rect 23714 14176 24034 15200
rect 23714 14112 23722 14176
rect 23786 14112 23802 14176
rect 23866 14112 23882 14176
rect 23946 14112 23962 14176
rect 24026 14112 24034 14176
rect 23714 13088 24034 14112
rect 23714 13024 23722 13088
rect 23786 13024 23802 13088
rect 23866 13024 23882 13088
rect 23946 13024 23962 13088
rect 24026 13024 24034 13088
rect 23714 12000 24034 13024
rect 23714 11936 23722 12000
rect 23786 11936 23802 12000
rect 23866 11936 23882 12000
rect 23946 11936 23962 12000
rect 24026 11936 24034 12000
rect 23714 10912 24034 11936
rect 23714 10848 23722 10912
rect 23786 10848 23802 10912
rect 23866 10848 23882 10912
rect 23946 10848 23962 10912
rect 24026 10848 24034 10912
rect 23714 9824 24034 10848
rect 23714 9760 23722 9824
rect 23786 9760 23802 9824
rect 23866 9760 23882 9824
rect 23946 9760 23962 9824
rect 24026 9760 24034 9824
rect 23714 8736 24034 9760
rect 23714 8672 23722 8736
rect 23786 8672 23802 8736
rect 23866 8672 23882 8736
rect 23946 8672 23962 8736
rect 24026 8672 24034 8736
rect 23714 7648 24034 8672
rect 23714 7584 23722 7648
rect 23786 7584 23802 7648
rect 23866 7584 23882 7648
rect 23946 7584 23962 7648
rect 24026 7584 24034 7648
rect 23714 6779 24034 7584
rect 23714 6560 23756 6779
rect 23992 6560 24034 6779
rect 23714 6496 23722 6560
rect 23786 6496 23802 6543
rect 23866 6496 23882 6543
rect 23946 6496 23962 6543
rect 24026 6496 24034 6560
rect 23714 5472 24034 6496
rect 23714 5408 23722 5472
rect 23786 5408 23802 5472
rect 23866 5408 23882 5472
rect 23946 5408 23962 5472
rect 24026 5408 24034 5472
rect 23714 4384 24034 5408
rect 23714 4320 23722 4384
rect 23786 4320 23802 4384
rect 23866 4320 23882 4384
rect 23946 4320 23962 4384
rect 24026 4320 24034 4384
rect 23714 3296 24034 4320
rect 26374 4045 26434 23427
rect 26371 4044 26437 4045
rect 26371 3980 26372 4044
rect 26436 3980 26437 4044
rect 26371 3979 26437 3980
rect 23714 3232 23722 3296
rect 23786 3232 23802 3296
rect 23866 3232 23882 3296
rect 23946 3232 23962 3296
rect 24026 3232 24034 3296
rect 23714 2208 24034 3232
rect 23714 2144 23722 2208
rect 23786 2144 23802 2208
rect 23866 2144 23882 2208
rect 23946 2144 23962 2208
rect 24026 2144 24034 2208
rect 23714 2128 24034 2144
<< via4 >>
rect 5540 24676 5776 24912
rect 10094 20160 10330 20379
rect 10094 20143 10124 20160
rect 10124 20143 10140 20160
rect 10140 20143 10204 20160
rect 10204 20143 10220 20160
rect 10220 20143 10284 20160
rect 10284 20143 10300 20160
rect 10300 20143 10330 20160
rect 5540 15610 5776 15846
rect 14648 24676 14884 24912
rect 10094 11076 10330 11312
rect 14648 15610 14884 15846
rect 5540 6560 5776 6779
rect 5540 6543 5570 6560
rect 5570 6543 5586 6560
rect 5586 6543 5650 6560
rect 5650 6543 5666 6560
rect 5666 6543 5730 6560
rect 5730 6543 5746 6560
rect 5746 6543 5776 6560
rect 14648 6560 14884 6779
rect 14648 6543 14678 6560
rect 14678 6543 14694 6560
rect 14694 6543 14758 6560
rect 14758 6543 14774 6560
rect 14774 6543 14838 6560
rect 14838 6543 14854 6560
rect 14854 6543 14884 6560
rect 19202 20160 19438 20379
rect 19202 20143 19232 20160
rect 19232 20143 19248 20160
rect 19248 20143 19312 20160
rect 19312 20143 19328 20160
rect 19328 20143 19392 20160
rect 19392 20143 19408 20160
rect 19408 20143 19438 20160
rect 19202 11076 19438 11312
rect 23756 24676 23992 24912
rect 23756 15610 23992 15846
rect 23756 6560 23992 6779
rect 23756 6543 23786 6560
rect 23786 6543 23802 6560
rect 23802 6543 23866 6560
rect 23866 6543 23882 6560
rect 23882 6543 23946 6560
rect 23946 6543 23962 6560
rect 23962 6543 23992 6560
<< metal5 >>
rect 1104 24912 28428 24955
rect 1104 24676 5540 24912
rect 5776 24676 14648 24912
rect 14884 24676 23756 24912
rect 23992 24676 28428 24912
rect 1104 24634 28428 24676
rect 1104 20379 28428 20421
rect 1104 20143 10094 20379
rect 10330 20143 19202 20379
rect 19438 20143 28428 20379
rect 1104 20101 28428 20143
rect 1104 15846 28428 15888
rect 1104 15610 5540 15846
rect 5776 15610 14648 15846
rect 14884 15610 23756 15846
rect 23992 15610 28428 15846
rect 1104 15568 28428 15610
rect 1104 11312 28428 11355
rect 1104 11076 10094 11312
rect 10330 11076 19202 11312
rect 19438 11076 28428 11312
rect 1104 11034 28428 11076
rect 1104 6779 28428 6821
rect 1104 6543 5540 6779
rect 5776 6543 14648 6779
rect 14884 6543 23756 6779
rect 23992 6543 28428 6779
rect 1104 6501 28428 6543
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1618216021
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618216021
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 1618216021
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1618216021
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1618216021
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1618216021
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11
timestamp 1618216021
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1618216021
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1033_
timestamp 1618216021
transform 1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1618216021
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17
timestamp 1618216021
transform 1 0 2668 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1618216021
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1037_
timestamp 1618216021
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1618216021
transform 1 0 3128 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1618216021
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1618216021
transform 1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1618216021
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1618216021
transform 1 0 4232 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1618216021
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1618216021
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1618216021
transform 1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1618216021
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1618216021
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1618216021
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1618216021
transform 1 0 4600 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1618216021
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1618216021
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1618216021
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1618216021
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1618216021
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1618216021
transform 1 0 6900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1618216021
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1618216021
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1618216021
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62
timestamp 1618216021
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_45
timestamp 1618216021
transform 1 0 5244 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1017_
timestamp 1618216021
transform 1 0 8004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1618216021
transform 1 0 7636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1618216021
transform 1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1618216021
transform 1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_66
timestamp 1618216021
transform 1 0 7176 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_74
timestamp 1618216021
transform 1 0 7912 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1618216021
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1618216021
transform 1 0 8372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1618216021
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1618216021
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1618216021
transform 1 0 8740 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1042_
timestamp 1618216021
transform 1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1618216021
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1618216021
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1618216021
transform 1 0 10856 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1618216021
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1618216021
transform 1 0 9936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1618216021
transform 1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_99
timestamp 1618216021
transform 1 0 10212 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1618216021
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1618216021
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1618216021
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1618216021
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1618216021
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1618216021
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_115
timestamp 1618216021
transform 1 0 11684 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1618216021
transform 1 0 12236 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_0_128
timestamp 1618216021
transform 1 0 12880 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1618216021
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1618216021
transform 1 0 12512 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1618216021
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136
timestamp 1618216021
transform 1 0 13616 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1618216021
transform 1 0 13984 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1618216021
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1618216021
transform 1 0 14352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1618216021
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1618216021
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1618216021
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1618216021
transform 1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1038_
timestamp 1618216021
transform 1 0 15088 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1005_
timestamp 1618216021
transform 1 0 15824 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_0_154
timestamp 1618216021
transform 1 0 15272 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1618216021
transform 1 0 15456 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1006_
timestamp 1618216021
transform 1 0 16008 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1618216021
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1618216021
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1618216021
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1618216021
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1618216021
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1618216021
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0939_
timestamp 1618216021
transform 1 0 18768 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1618216021
transform 1 0 17296 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1618216021
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1618216021
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_183
timestamp 1618216021
transform 1 0 17940 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp 1618216021
transform 1 0 18676 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_192
timestamp 1618216021
transform 1 0 18768 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1618216021
transform 1 0 19320 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1618216021
transform 1 0 20608 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1618216021
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1618216021
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1618216021
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_204
timestamp 1618216021
transform 1 0 19872 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1618216021
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0937_
timestamp 1618216021
transform 1 0 22908 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1618216021
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1618216021
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1618216021
transform 1 0 22540 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1618216021
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1618216021
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_222
timestamp 1618216021
transform 1 0 21528 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1618216021
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1618216021
transform 1 0 22908 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1618216021
transform 1 0 23460 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1618216021
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1618216021
transform 1 0 23920 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1618216021
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_252
timestamp 1618216021
transform 1 0 24288 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_260
timestamp 1618216021
transform 1 0 25024 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1618216021
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_259
timestamp 1618216021
transform 1 0 24932 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1618216021
transform 1 0 25576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1618216021
transform 1 0 25852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1618216021
transform 1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_267
timestamp 1618216021
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1618216021
transform 1 0 26312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_273
timestamp 1618216021
transform 1 0 26220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1618216021
transform 1 0 26588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_278
timestamp 1618216021
transform 1 0 26680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1618216021
transform 1 0 26956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1618216021
transform 1 0 27048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618216021
transform -1 0 28428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618216021
transform -1 0 28428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1618216021
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1618216021
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1618216021
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_291
timestamp 1618216021
transform 1 0 27876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_286
timestamp 1618216021
transform 1 0 27416 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1035_
timestamp 1618216021
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618216021
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1618216021
transform 1 0 2852 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1618216021
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1618216021
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1618216021
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1618216021
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1618216021
transform 1 0 3128 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_28
timestamp 1618216021
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1618216021
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_42
timestamp 1618216021
transform 1 0 4968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1618216021
transform 1 0 5520 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_64
timestamp 1618216021
transform 1 0 6992 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1618216021
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1618216021
transform 1 0 8372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1618216021
transform 1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1618216021
transform 1 0 8004 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1618216021
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_87
timestamp 1618216021
transform 1 0 9108 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0955_
timestamp 1618216021
transform 1 0 9936 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1618216021
transform 1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_95
timestamp 1618216021
transform 1 0 9844 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1618216021
transform 1 0 10580 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0902_
timestamp 1618216021
transform 1 0 12788 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1618216021
transform 1 0 12420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1618216021
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output150
timestamp 1618216021
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_134
timestamp 1618216021
transform 1 0 13432 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1618216021
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1618216021
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_148
timestamp 1618216021
transform 1 0 14720 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1618216021
transform 1 0 15548 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1618216021
transform 1 0 15180 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1618216021
transform 1 0 17020 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1618216021
transform 1 0 18124 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1618216021
transform 1 0 17388 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1618216021
transform 1 0 18768 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1618216021
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp 1618216021
transform 1 0 18032 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_188
timestamp 1618216021
transform 1 0 18400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_196
timestamp 1618216021
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1618216021
transform 1 0 19964 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0936_
timestamp 1618216021
transform 1 0 20608 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1618216021
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1618216021
transform 1 0 19596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1618216021
transform 1 0 20240 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1618216021
transform 1 0 21620 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1618216021
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1618216021
transform 1 0 23092 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1002_
timestamp 1618216021
transform 1 0 23460 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1618216021
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_250
timestamp 1618216021
transform 1 0 24104 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_256
timestamp 1618216021
transform 1 0 24656 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1618216021
transform 1 0 24840 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1015_
timestamp 1618216021
transform 1 0 26956 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1618216021
transform 1 0 26220 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1618216021
transform 1 0 25484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_264
timestamp 1618216021
transform 1 0 25392 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_269
timestamp 1618216021
transform 1 0 25852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1618216021
transform 1 0 26588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618216021
transform -1 0 28428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_285
timestamp 1618216021
transform 1 0 27324 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_293
timestamp 1618216021
transform 1 0 28060 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618216021
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1618216021
transform 1 0 2484 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1618216021
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1618216021
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1618216021
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1618216021
transform 1 0 2760 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1618216021
transform 1 0 4324 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1618216021
transform 1 0 3128 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_25
timestamp 1618216021
transform 1 0 3404 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1618216021
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1618216021
transform 1 0 4968 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0907_
timestamp 1618216021
transform 1 0 5336 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1618216021
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1618216021
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1618216021
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1618216021
transform 1 0 8924 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1618216021
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_82
timestamp 1618216021
transform 1 0 8648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output160
timestamp 1618216021
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1618216021
transform 1 0 10396 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_109
timestamp 1618216021
transform 1 0 11132 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1618216021
transform 1 0 12052 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1618216021
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1618216021
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1618216021
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1618216021
transform 1 0 13892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1618216021
transform 1 0 14536 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1618216021
transform 1 0 13524 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1618216021
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1618216021
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1618216021
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1618216021
transform 1 0 15180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1618216021
transform 1 0 16100 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_156
timestamp 1618216021
transform 1 0 15456 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp 1618216021
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1618216021
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1618216021
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1618216021
transform 1 0 17296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0999_
timestamp 1618216021
transform 1 0 17940 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1618216021
transform 1 0 18952 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1618216021
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1618216021
transform 1 0 18584 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1618216021
transform 1 0 21160 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_210
timestamp 1618216021
transform 1 0 20424 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1618216021
transform 1 0 22540 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1618216021
transform 1 0 23184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1618216021
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_221
timestamp 1618216021
transform 1 0 21436 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_227
timestamp 1618216021
transform 1 0 21988 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1618216021
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_236
timestamp 1618216021
transform 1 0 22816 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1618216021
transform 1 0 23828 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1618216021
transform 1 0 24840 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1618216021
transform 1 0 23460 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_250
timestamp 1618216021
transform 1 0 24104 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_261
timestamp 1618216021
transform 1 0 25116 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1618216021
transform 1 0 25944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output153
timestamp 1618216021
transform 1 0 26588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_269
timestamp 1618216021
transform 1 0 25852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_273
timestamp 1618216021
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1618216021
transform 1 0 26956 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618216021
transform -1 0 28428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1618216021
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_286
timestamp 1618216021
transform 1 0 27416 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0911_
timestamp 1618216021
transform 1 0 2300 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618216021
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1618216021
transform 1 0 1564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1618216021
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1618216021
transform 1 0 1932 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1618216021
transform 1 0 2944 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1618216021
transform 1 0 4784 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1618216021
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1618216021
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_30
timestamp 1618216021
transform 1 0 3864 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_38
timestamp 1618216021
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1618216021
transform 1 0 6716 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1618216021
transform 1 0 6256 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1618216021
transform 1 0 6624 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_64
timestamp 1618216021
transform 1 0 6992 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1618216021
transform 1 0 8372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1618216021
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_76
timestamp 1618216021
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1618216021
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1618216021
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1618216021
transform 1 0 9568 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1618216021
transform 1 0 11040 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1618216021
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_99
timestamp 1618216021
transform 1 0 10212 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_107
timestamp 1618216021
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0953_
timestamp 1618216021
transform 1 0 12880 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1618216021
transform 1 0 12512 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp 1618216021
transform 1 0 14720 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1618216021
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1618216021
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1618216021
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1618216021
transform 1 0 16928 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_164
timestamp 1618216021
transform 1 0 16192 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1618216021
transform 1 0 17664 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_176
timestamp 1618216021
transform 1 0 17296 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1618216021
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0942_
timestamp 1618216021
transform 1 0 19964 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1618216021
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1618216021
transform 1 0 20976 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1618216021
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_212
timestamp 1618216021
transform 1 0 20608 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1618216021
transform 1 0 22816 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1618216021
transform 1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1618216021
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_226
timestamp 1618216021
transform 1 0 21896 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_234
timestamp 1618216021
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1618216021
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1618216021
transform 1 0 25208 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_252
timestamp 1618216021
transform 1 0 24288 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_256
timestamp 1618216021
transform 1 0 24656 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1618216021
transform 1 0 24840 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1618216021
transform 1 0 26772 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1618216021
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_265
timestamp 1618216021
transform 1 0 25484 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_271
timestamp 1618216021
transform 1 0 26036 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1618216021
transform 1 0 26404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1618216021
transform 1 0 27048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618216021
transform -1 0 28428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1618216021
transform 1 0 27416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_290
timestamp 1618216021
transform 1 0 27784 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1618216021
transform 1 0 2116 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1618216021
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1618216021
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1618216021
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_10
timestamp 1618216021
transform 1 0 2024 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1618216021
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1618216021
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1618216021
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1618216021
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1618216021
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_58
timestamp 1618216021
transform 1 0 6440 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_64
timestamp 1618216021
transform 1 0 6992 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1618216021
transform 1 0 7728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1618216021
transform 1 0 8372 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1618216021
transform 1 0 7360 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_75
timestamp 1618216021
transform 1 0 8004 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0808_
timestamp 1618216021
transform 1 0 10212 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1618216021
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1618216021
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0806_
timestamp 1618216021
transform 1 0 12052 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1618216021
transform 1 0 13064 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1618216021
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1618216021
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1618216021
transform 1 0 12696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1618216021
transform 1 0 14996 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_147
timestamp 1618216021
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0997_
timestamp 1618216021
transform 1 0 15824 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1618216021
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_154
timestamp 1618216021
transform 1 0 15272 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1618216021
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1618216021
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0941_
timestamp 1618216021
transform 1 0 17296 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0998_
timestamp 1618216021
transform 1 0 18032 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1618216021
transform 1 0 19044 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_180
timestamp 1618216021
transform 1 0 17664 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1618216021
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_211
timestamp 1618216021
transform 1 0 20516 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1618216021
transform 1 0 21436 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1004_
timestamp 1618216021
transform 1 0 22632 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1618216021
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_219
timestamp 1618216021
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_224
timestamp 1618216021
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1618216021
transform 1 0 22172 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1618216021
transform 1 0 22540 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1618216021
transform 1 0 23736 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_241
timestamp 1618216021
transform 1 0 23276 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_245
timestamp 1618216021
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1618216021
transform 1 0 25208 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1618216021
transform 1 0 26680 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_274
timestamp 1618216021
transform 1 0 26312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1618216021
transform 1 0 26956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1618216021
transform -1 0 28428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1618216021
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_286
timestamp 1618216021
transform 1 0 27416 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1618216021
transform 1 0 2852 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1618216021
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1618216021
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1618216021
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1618216021
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1618216021
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_6
timestamp 1618216021
transform 1 0 1656 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_18
timestamp 1618216021
transform 1 0 2760 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1618216021
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0906_
timestamp 1618216021
transform 1 0 4692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1618216021
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1618216021
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1618216021
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_37
timestamp 1618216021
transform 1 0 4508 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1618216021
transform 1 0 4324 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1618216021
transform 1 0 5060 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0899_
timestamp 1618216021
transform 1 0 5428 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1618216021
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_49
timestamp 1618216021
transform 1 0 5612 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1618216021
transform 1 0 6716 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_65
timestamp 1618216021
transform 1 0 7084 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1618216021
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1618216021
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _0562_
timestamp 1618216021
transform 1 0 7912 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0563_
timestamp 1618216021
transform 1 0 8924 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 1618216021
transform 1 0 7176 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1618216021
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_82
timestamp 1618216021
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1618216021
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1618216021
transform 1 0 7544 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1618216021
transform 1 0 8556 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1618216021
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0564_
timestamp 1618216021
transform 1 0 9476 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 1618216021
transform 1 0 10120 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1618216021
transform 1 0 10764 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_109
timestamp 1618216021
transform 1 0 11132 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_92
timestamp 1618216021
transform 1 0 9568 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1618216021
transform 1 0 10672 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0547_
timestamp 1618216021
transform 1 0 12788 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0548_
timestamp 1618216021
transform 1 0 12604 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0854_
timestamp 1618216021
transform 1 0 11224 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1618216021
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_117
timestamp 1618216021
transform 1 0 11868 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1618216021
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1618216021
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_115
timestamp 1618216021
transform 1 0 11684 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1618216021
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1618216021
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0549_
timestamp 1618216021
transform 1 0 13984 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1618216021
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_134
timestamp 1618216021
transform 1 0 13432 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1618216021
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1618216021
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_151
timestamp 1618216021
transform 1 0 14996 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_132
timestamp 1618216021
transform 1 0 13248 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_147
timestamp 1618216021
transform 1 0 14628 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0943_
timestamp 1618216021
transform 1 0 15824 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1618216021
transform 1 0 15456 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1618216021
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1618216021
transform 1 0 15180 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_155
timestamp 1618216021
transform 1 0 15364 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_172
timestamp 1618216021
transform 1 0 16928 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1618216021
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1618216021
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_172
timestamp 1618216021
transform 1 0 16928 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1618216021
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0940_
timestamp 1618216021
transform 1 0 17480 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_7_182
timestamp 1618216021
transform 1 0 17848 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0933_
timestamp 1618216021
transform 1 0 19044 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0934_
timestamp 1618216021
transform 1 0 18768 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1001_
timestamp 1618216021
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_188
timestamp 1618216021
transform 1 0 18400 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1618216021
transform 1 0 19136 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_190
timestamp 1618216021
transform 1 0 18584 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_194
timestamp 1618216021
transform 1 0 18952 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _0745_
timestamp 1618216021
transform 1 0 21068 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0938_
timestamp 1618216021
transform 1 0 20516 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1618216021
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1618216021
transform 1 0 19964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1618216021
transform 1 0 19596 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_208
timestamp 1618216021
transform 1 0 20240 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_216
timestamp 1618216021
transform 1 0 20976 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_199
timestamp 1618216021
transform 1 0 19412 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_218
timestamp 1618216021
transform 1 0 21160 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0755_
timestamp 1618216021
transform 1 0 23092 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0762_
timestamp 1618216021
transform 1 0 22540 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1618216021
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_223
timestamp 1618216021
transform 1 0 21620 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_231
timestamp 1618216021
transform 1 0 22356 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_239
timestamp 1618216021
transform 1 0 23092 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_226
timestamp 1618216021
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_229
timestamp 1618216021
transform 1 0 22172 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_237
timestamp 1618216021
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _0754_
timestamp 1618216021
transform 1 0 24288 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1003_
timestamp 1618216021
transform 1 0 23460 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1618216021
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_250
timestamp 1618216021
transform 1 0 24104 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_256
timestamp 1618216021
transform 1 0 24656 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1618216021
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1618216021
transform 1 0 23920 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_258
timestamp 1618216021
transform 1 0 24840 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1618216021
transform 1 0 26588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_270
timestamp 1618216021
transform 1 0 25944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1618216021
transform 1 0 27048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_270
timestamp 1618216021
transform 1 0 25944 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1618216021
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1618216021
transform 1 0 26956 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1618216021
transform -1 0 28428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1618216021
transform -1 0 28428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1618216021
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1618216021
transform 1 0 27416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_290
timestamp 1618216021
transform 1 0 27784 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_286
timestamp 1618216021
transform 1 0 27416 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1618216021
transform 1 0 1748 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1618216021
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1618216021
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0909_
timestamp 1618216021
transform 1 0 4232 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1618216021
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_23
timestamp 1618216021
transform 1 0 3220 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1618216021
transform 1 0 3864 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1618216021
transform 1 0 4876 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1618216021
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0905_
timestamp 1618216021
transform 1 0 5428 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1618216021
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_58
timestamp 1618216021
transform 1 0 6440 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0569_
timestamp 1618216021
transform 1 0 7176 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1618216021
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_73
timestamp 1618216021
transform 1 0 7820 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1618216021
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1618216021
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0855_
timestamp 1618216021
transform 1 0 10856 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_8_99
timestamp 1618216021
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp 1618216021
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1618216021
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_113
timestamp 1618216021
transform 1 0 11500 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_119
timestamp 1618216021
transform 1 0 12052 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1618216021
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1618216021
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1618216021
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1618216021
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1618216021
transform 1 0 15732 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp 1618216021
transform 1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1618216021
transform 1 0 18032 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1618216021
transform 1 0 18676 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_175
timestamp 1618216021
transform 1 0 17204 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1618216021
transform 1 0 17940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_187
timestamp 1618216021
transform 1 0 18308 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_194
timestamp 1618216021
transform 1 0 18952 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1618216021
transform 1 0 20148 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1618216021
transform 1 0 20792 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1618216021
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_201
timestamp 1618216021
transform 1 0 19596 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1618216021
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1618216021
transform 1 0 22632 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1618216021
transform 1 0 22264 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0988_
timestamp 1618216021
transform 1 0 25208 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1618216021
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_250
timestamp 1618216021
transform 1 0 24104 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_256
timestamp 1618216021
transform 1 0 24656 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1618216021
transform 1 0 24840 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1063_
timestamp 1618216021
transform 1 0 26220 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_8_269
timestamp 1618216021
transform 1 0 25852 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1618216021
transform -1 0 28428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_290
timestamp 1618216021
transform 1 0 27784 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0908_
timestamp 1618216021
transform 1 0 2116 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1618216021
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1618216021
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1618216021
transform 1 0 1748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_18
timestamp 1618216021
transform 1 0 2760 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0586_
timestamp 1618216021
transform 1 0 3496 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1618216021
transform 1 0 4416 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1618216021
transform 1 0 4048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0578_
timestamp 1618216021
transform 1 0 6808 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1618216021
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1618216021
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_56
timestamp 1618216021
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_58
timestamp 1618216021
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1618216021
transform 1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1618216021
transform 1 0 7452 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_76
timestamp 1618216021
transform 1 0 8096 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _0555_
timestamp 1618216021
transform 1 0 10580 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_88
timestamp 1618216021
transform 1 0 9200 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_100
timestamp 1618216021
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1618216021
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1618216021
transform 1 0 12696 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1618216021
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1618216021
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1618216021
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1618216021
transform 1 0 12328 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_129
timestamp 1618216021
transform 1 0 12972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1618216021
transform 1 0 14076 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1618216021
transform 1 0 16192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1618216021
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1618216021
transform 1 0 15180 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_161
timestamp 1618216021
transform 1 0 15916 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1618216021
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_172
timestamp 1618216021
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1061_
timestamp 1618216021
transform 1 0 17664 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__or2b_1  _0736_
timestamp 1618216021
transform 1 0 19596 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0935_
timestamp 1618216021
transform 1 0 21068 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1618216021
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_207
timestamp 1618216021
transform 1 0 20148 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1618216021
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _0746_
timestamp 1618216021
transform 1 0 22540 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1618216021
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_224
timestamp 1618216021
transform 1 0 21712 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1618216021
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0987_
timestamp 1618216021
transform 1 0 23828 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1064_
timestamp 1618216021
transform 1 0 24840 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_9_242
timestamp 1618216021
transform 1 0 23368 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_246
timestamp 1618216021
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_254
timestamp 1618216021
transform 1 0 24472 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_275
timestamp 1618216021
transform 1 0 26404 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1618216021
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1618216021
transform -1 0 28428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1618216021
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_286
timestamp 1618216021
transform 1 0 27416 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1032_
timestamp 1618216021
transform 1 0 2116 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1618216021
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1618216021
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1618216021
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_10
timestamp 1618216021
transform 1 0 2024 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1618216021
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0860_
timestamp 1618216021
transform 1 0 4416 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1618216021
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1618216021
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_30
timestamp 1618216021
transform 1 0 3864 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_43
timestamp 1618216021
transform 1 0 5060 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1618216021
transform 1 0 5428 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1618216021
transform 1 0 6900 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0859_
timestamp 1618216021
transform 1 0 7268 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1618216021
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1618216021
transform 1 0 7912 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_87
timestamp 1618216021
transform 1 0 9108 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1618216021
transform 1 0 10488 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_i_clk
timestamp 1618216021
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_98
timestamp 1618216021
transform 1 0 10120 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1618216021
transform 1 0 12328 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1618216021
transform 1 0 11960 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp 1618216021
transform 1 0 14720 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1618216021
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_138
timestamp 1618216021
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1618216021
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1618216021
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0728_
timestamp 1618216021
transform 1 0 16560 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1618216021
transform 1 0 16192 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1618216021
transform 1 0 17112 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1618216021
transform 1 0 18492 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0990_
timestamp 1618216021
transform 1 0 17480 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1618216021
transform 1 0 18124 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_196
timestamp 1618216021
transform 1 0 19136 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0737_
timestamp 1618216021
transform 1 0 20424 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1618216021
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_201
timestamp 1618216021
transform 1 0 19596 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1618216021
transform 1 0 20332 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1618216021
transform 1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0763_
timestamp 1618216021
transform 1 0 22632 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1618216021
transform 1 0 21252 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_226
timestamp 1618216021
transform 1 0 21896 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1618216021
transform 1 0 25208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1618216021
transform 1 0 24104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1618216021
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_243
timestamp 1618216021
transform 1 0 23460 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_249
timestamp 1618216021
transform 1 0 24012 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1618216021
transform 1 0 24380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1618216021
transform 1 0 24840 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1062_
timestamp 1618216021
transform 1 0 25944 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1618216021
transform 1 0 25484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_269
timestamp 1618216021
transform 1 0 25852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1618216021
transform -1 0 28428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_287
timestamp 1618216021
transform 1 0 27508 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1618216021
transform 1 0 28060 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0962_
timestamp 1618216021
transform 1 0 2300 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1618216021
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1618216021
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1618216021
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_20
timestamp 1618216021
transform 1 0 2944 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0602_
timestamp 1618216021
transform 1 0 3864 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1618216021
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_36
timestamp 1618216021
transform 1 0 4416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1618216021
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1618216021
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1618216021
transform 1 0 5520 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1618216021
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_58
timestamp 1618216021
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_65
timestamp 1618216021
transform 1 0 7084 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1618216021
transform 1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 1618216021
transform 1 0 8188 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_69
timestamp 1618216021
transform 1 0 7452 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1618216021
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0570_
timestamp 1618216021
transform 1 0 10028 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1618216021
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_109
timestamp 1618216021
transform 1 0 11132 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1618216021
transform 1 0 12052 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1618216021
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1618216021
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1618216021
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_126
timestamp 1618216021
transform 1 0 12696 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0571_
timestamp 1618216021
transform 1 0 13340 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 1618216021
transform 1 0 14352 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_132
timestamp 1618216021
transform 1 0 13248 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1618216021
transform 1 0 13984 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1618216021
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1618216021
transform 1 0 15824 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_168
timestamp 1618216021
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1618216021
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0727_
timestamp 1618216021
transform 1 0 17296 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1618216021
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1065_
timestamp 1618216021
transform 1 0 18768 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1618216021
transform 1 0 17664 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1618216021
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1618216021
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1618216021
transform 1 0 20700 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1618216021
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_216
timestamp 1618216021
transform 1 0 20976 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1618216021
transform 1 0 22724 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1618216021
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_i_clk
timestamp 1618216021
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_223
timestamp 1618216021
transform 1 0 21620 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_227
timestamp 1618216021
transform 1 0 21988 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_229
timestamp 1618216021
transform 1 0 22172 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_238
timestamp 1618216021
transform 1 0 23000 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1618216021
transform 1 0 24564 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_i_clk
timestamp 1618216021
transform 1 0 23920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_246
timestamp 1618216021
transform 1 0 23736 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1618216021
transform 1 0 24196 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_262
timestamp 1618216021
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0989_
timestamp 1618216021
transform 1 0 25576 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1618216021
transform 1 0 26680 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_273
timestamp 1618216021
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_277
timestamp 1618216021
transform 1 0 26588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1618216021
transform 1 0 26956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1618216021
transform -1 0 28428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1618216021
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_286
timestamp 1618216021
transform 1 0 27416 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0959_
timestamp 1618216021
transform 1 0 2116 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1618216021
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1618216021
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1618216021
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_10
timestamp 1618216021
transform 1 0 2024 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_18
timestamp 1618216021
transform 1 0 2760 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1618216021
transform 1 0 3128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1618216021
transform 1 0 5060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1618216021
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1618216021
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_25
timestamp 1618216021
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_30
timestamp 1618216021
transform 1 0 3864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_34
timestamp 1618216021
transform 1 0 4232 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1618216021
transform 1 0 4600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_42
timestamp 1618216021
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1618216021
transform 1 0 6348 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_i_clk
timestamp 1618216021
transform 1 0 5704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1618216021
transform 1 0 5336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 1618216021
transform 1 0 5980 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_64
timestamp 1618216021
transform 1 0 6992 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_2  _0579_
timestamp 1618216021
transform 1 0 7544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1618216021
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_82
timestamp 1618216021
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1618216021
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0556_
timestamp 1618216021
transform 1 0 10856 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0557_
timestamp 1618216021
transform 1 0 9476 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_98
timestamp 1618216021
transform 1 0 10120 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0544_
timestamp 1618216021
transform 1 0 12604 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_118
timestamp 1618216021
transform 1 0 11960 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_124
timestamp 1618216021
transform 1 0 12512 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1618216021
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0541_
timestamp 1618216021
transform 1 0 13340 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0580_
timestamp 1618216021
transform 1 0 14720 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1618216021
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_137
timestamp 1618216021
transform 1 0 13708 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1618216021
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0895_
timestamp 1618216021
transform 1 0 16560 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_155
timestamp 1618216021
transform 1 0 15364 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1618216021
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_172
timestamp 1618216021
transform 1 0 16928 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0984_
timestamp 1618216021
transform 1 0 17572 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0985_
timestamp 1618216021
transform 1 0 18308 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_178
timestamp 1618216021
transform 1 0 17480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1618216021
transform 1 0 17940 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_191
timestamp 1618216021
transform 1 0 18676 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0891_
timestamp 1618216021
transform 1 0 19964 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1618216021
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1618216021
transform 1 0 19412 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1618216021
transform 1 0 19596 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_212
timestamp 1618216021
transform 1 0 20608 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0889_
timestamp 1618216021
transform 1 0 22724 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_224
timestamp 1618216021
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_232
timestamp 1618216021
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1618216021
transform 1 0 24104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0841_
timestamp 1618216021
transform 1 0 25208 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1618216021
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_242
timestamp 1618216021
transform 1 0 23368 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1618216021
transform 1 0 24380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1618216021
transform 1 0 24840 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1618216021
transform 1 0 26772 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_269
timestamp 1618216021
transform 1 0 25852 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_277
timestamp 1618216021
transform 1 0 26588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_282
timestamp 1618216021
transform 1 0 27048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1618216021
transform -1 0 28428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1618216021
transform 1 0 27416 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1618216021
transform 1 0 27784 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1081_
timestamp 1618216021
transform 1 0 2024 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1618216021
transform 1 0 1472 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1618216021
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1618216021
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1618216021
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1618216021
transform 1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1618216021
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1618216021
transform 1 0 2944 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0815_
timestamp 1618216021
transform 1 0 3956 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1618216021
transform 1 0 4232 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1618216021
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1618216021
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_38
timestamp 1618216021
transform 1 0 4600 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_28
timestamp 1618216021
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_30
timestamp 1618216021
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0812_
timestamp 1618216021
transform 1 0 5336 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1618216021
transform 1 0 6072 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1618216021
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1618216021
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_53
timestamp 1618216021
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_58
timestamp 1618216021
transform 1 0 6440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_50
timestamp 1618216021
transform 1 0 5704 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1618216021
transform 1 0 8648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1618216021
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1618216021
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1618216021
transform 1 0 8924 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1618216021
transform 1 0 7544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1618216021
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1618216021
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0536_
timestamp 1618216021
transform 1 0 9476 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1618216021
transform 1 0 9292 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_i_clk
timestamp 1618216021
transform 1 0 10028 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_92
timestamp 1618216021
transform 1 0 9568 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_96
timestamp 1618216021
transform 1 0 9936 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_98
timestamp 1618216021
transform 1 0 10120 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1618216021
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1618216021
transform 1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_100
timestamp 1618216021
transform 1 0 10304 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_106
timestamp 1618216021
transform 1 0 10856 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1618216021
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0954_
timestamp 1618216021
transform 1 0 11868 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1087_
timestamp 1618216021
transform 1 0 12420 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1618216021
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1618216021
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_115
timestamp 1618216021
transform 1 0 11684 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_124
timestamp 1618216021
transform 1 0 12512 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0537_
timestamp 1618216021
transform 1 0 14352 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1618216021
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1618216021
transform 1 0 13984 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_148
timestamp 1618216021
transform 1 0 14720 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_136
timestamp 1618216021
transform 1 0 13616 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1618216021
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1618216021
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1618216021
transform 1 0 16192 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1618216021
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1618216021
transform 1 0 15824 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_168
timestamp 1618216021
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_172
timestamp 1618216021
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_156
timestamp 1618216021
transform 1 0 15456 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0773_
timestamp 1618216021
transform 1 0 18124 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _0775_
timestamp 1618216021
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 1618216021
transform 1 0 17296 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_185
timestamp 1618216021
transform 1 0 18124 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1618216021
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 1618216021
transform 1 0 18032 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1618216021
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1618216021
transform 1 0 21160 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0843_
timestamp 1618216021
transform 1 0 20148 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1618216021
transform 1 0 19964 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1618216021
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1618216021
transform 1 0 19780 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_214
timestamp 1618216021
transform 1 0 20792 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1618216021
transform 1 0 19596 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0764_
timestamp 1618216021
transform 1 0 22908 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1618216021
transform 1 0 22264 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1618216021
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_221
timestamp 1618216021
transform 1 0 21436 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_227
timestamp 1618216021
transform 1 0 21988 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_229
timestamp 1618216021
transform 1 0 22172 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_221
timestamp 1618216021
transform 1 0 21436 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_229
timestamp 1618216021
transform 1 0 22172 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1618216021
transform 1 0 24104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1618216021
transform 1 0 24840 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1618216021
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1618216021
transform 1 0 24012 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_257
timestamp 1618216021
transform 1 0 24748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_246
timestamp 1618216021
transform 1 0 23736 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1618216021
transform 1 0 24380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1618216021
transform 1 0 24840 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_262
timestamp 1618216021
transform 1 0 25208 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1618216021
transform 1 0 25300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1618216021
transform 1 0 26680 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_274
timestamp 1618216021
transform 1 0 26312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1618216021
transform 1 0 26956 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_279
timestamp 1618216021
transform 1 0 26772 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1618216021
transform -1 0 28428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1618216021
transform -1 0 28428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1618216021
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1618216021
transform 1 0 27416 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_286
timestamp 1618216021
transform 1 0 27416 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_285
timestamp 1618216021
transform 1 0 27324 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_290
timestamp 1618216021
transform 1 0 27784 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1618216021
transform 1 0 2668 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1618216021
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1618216021
transform 1 0 1748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1618216021
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_11
timestamp 1618216021
transform 1 0 2116 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0603_
timestamp 1618216021
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_33
timestamp 1618216021
transform 1 0 4140 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _0604_
timestamp 1618216021
transform 1 0 6808 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1618216021
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1618216021
transform 1 0 5520 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1618216021
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_58
timestamp 1618216021
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 1618216021
transform 1 0 8740 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1618216021
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0805_
timestamp 1618216021
transform 1 0 10580 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1618216021
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1618216021
transform 1 0 12052 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1618216021
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1618216021
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1618216021
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0511_
timestamp 1618216021
transform 1 0 13892 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp 1618216021
transform 1 0 14628 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1618216021
transform 1 0 13524 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_143
timestamp 1618216021
transform 1 0 14260 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1618216021
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1618216021
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1618216021
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0774_
timestamp 1618216021
transform 1 0 17848 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_180
timestamp 1618216021
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_191
timestamp 1618216021
transform 1 0 18676 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1618216021
transform 1 0 19596 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1618216021
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_217
timestamp 1618216021
transform 1 0 21068 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1618216021
transform 1 0 22724 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1618216021
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1618216021
transform 1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_229
timestamp 1618216021
transform 1 0 22172 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1618216021
transform 1 0 24840 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_251
timestamp 1618216021
transform 1 0 24196 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_257
timestamp 1618216021
transform 1 0 24748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1618216021
transform 1 0 25116 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp 1618216021
transform 1 0 25484 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1618216021
transform 1 0 26956 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1618216021
transform -1 0 28428 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1618216021
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_286
timestamp 1618216021
transform 1 0 27416 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1618216021
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1618216021
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1618216021
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0863_
timestamp 1618216021
transform 1 0 4232 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1618216021
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1618216021
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1618216021
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1618216021
transform 1 0 4876 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1618216021
transform 1 0 5704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_i_clk
timestamp 1618216021
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_49
timestamp 1618216021
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1618216021
transform 1 0 5980 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 1618216021
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o211ai_1  _0535_
timestamp 1618216021
transform 1 0 8096 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1618216021
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_66
timestamp 1618216021
transform 1 0 7176 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_74
timestamp 1618216021
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_82
timestamp 1618216021
transform 1 0 8648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_87
timestamp 1618216021
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1618216021
transform 1 0 10028 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_95
timestamp 1618216021
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0518_
timestamp 1618216021
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0804_
timestamp 1618216021
transform 1 0 11868 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_113
timestamp 1618216021
transform 1 0 11500 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_124
timestamp 1618216021
transform 1 0 12512 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1618216021
transform 1 0 13616 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1014_
timestamp 1618216021
transform 1 0 14720 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1618216021
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_132
timestamp 1618216021
transform 1 0 13248 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1618216021
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1618216021
transform 1 0 14352 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0572_
timestamp 1618216021
transform 1 0 15732 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0796_
timestamp 1618216021
transform 1 0 16744 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1618216021
transform 1 0 15364 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_163
timestamp 1618216021
transform 1 0 16100 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_169
timestamp 1618216021
transform 1 0 16652 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0517_
timestamp 1618216021
transform 1 0 18032 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1618216021
transform 1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_177
timestamp 1618216021
transform 1 0 17388 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1618216021
transform 1 0 17940 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_188
timestamp 1618216021
transform 1 0 18400 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_192
timestamp 1618216021
transform 1 0 18768 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_196
timestamp 1618216021
transform 1 0 19136 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0887_
timestamp 1618216021
transform 1 0 20516 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1618216021
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_201
timestamp 1618216021
transform 1 0 19596 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_209
timestamp 1618216021
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_218
timestamp 1618216021
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0890_
timestamp 1618216021
transform 1 0 22264 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1618216021
transform 1 0 22908 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0756_
timestamp 1618216021
transform 1 0 23276 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1618216021
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1618216021
transform 1 0 24380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1618216021
transform 1 0 24840 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_262
timestamp 1618216021
transform 1 0 25208 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0605_
timestamp 1618216021
transform 1 0 25300 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp 1618216021
transform 1 0 26312 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1618216021
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1618216021
transform -1 0 28428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_290
timestamp 1618216021
transform 1 0 27784 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1025_
timestamp 1618216021
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1618216021
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output152
timestamp 1618216021
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1618216021
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1618216021
transform 1 0 2484 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1618216021
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1618216021
transform 1 0 4140 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0813_
timestamp 1618216021
transform 1 0 3128 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1618216021
transform 1 0 3772 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_36
timestamp 1618216021
transform 1 0 4416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0809_
timestamp 1618216021
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1618216021
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_i_clk
timestamp 1618216021
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1618216021
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1618216021
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0583_
timestamp 1618216021
transform 1 0 8372 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_66
timestamp 1618216021
transform 1 0 7176 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_78
timestamp 1618216021
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1618216021
transform 1 0 8924 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1618216021
transform 1 0 9292 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_105
timestamp 1618216021
transform 1 0 10764 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0800_
timestamp 1618216021
transform 1 0 12052 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _1013_
timestamp 1618216021
transform 1 0 13156 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1618216021
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1618216021
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1618216021
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1618216021
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_143
timestamp 1618216021
transform 1 0 14260 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0894_
timestamp 1618216021
transform 1 0 15732 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1618216021
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1618216021
transform 1 0 15364 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_164
timestamp 1618216021
transform 1 0 16192 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_170
timestamp 1618216021
transform 1 0 16744 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_172
timestamp 1618216021
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1618216021
transform 1 0 17296 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1618216021
transform 1 0 18768 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_196
timestamp 1618216021
transform 1 0 19136 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0839_
timestamp 1618216021
transform 1 0 20608 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_i_clk
timestamp 1618216021
transform 1 0 19228 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_i_clk
timestamp 1618216021
transform 1 0 19872 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1618216021
transform 1 0 19504 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_207
timestamp 1618216021
transform 1 0 20148 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1618216021
transform 1 0 20516 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1618216021
transform 1 0 23184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1618216021
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_219
timestamp 1618216021
transform 1 0 21252 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_227
timestamp 1618216021
transform 1 0 21988 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_229
timestamp 1618216021
transform 1 0 22172 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_237
timestamp 1618216021
transform 1 0 22908 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1618216021
transform 1 0 24748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_i_clk
timestamp 1618216021
transform 1 0 23828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1618216021
transform 1 0 23460 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_250
timestamp 1618216021
transform 1 0 24104 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_256
timestamp 1618216021
transform 1 0 24656 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1618216021
transform 1 0 25024 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0613_
timestamp 1618216021
transform 1 0 26036 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_i_clk
timestamp 1618216021
transform 1 0 25392 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_267
timestamp 1618216021
transform 1 0 25668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_278
timestamp 1618216021
transform 1 0 26680 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1618216021
transform -1 0 28428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1618216021
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_284
timestamp 1618216021
transform 1 0 27232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_286
timestamp 1618216021
transform 1 0 27416 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1618216021
transform 1 0 1932 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1618216021
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1618216021
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0587_
timestamp 1618216021
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1618216021
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_25
timestamp 1618216021
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_30
timestamp 1618216021
transform 1 0 3864 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1618216021
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_2  _0588_
timestamp 1618216021
transform 1 0 5796 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0810_
timestamp 1618216021
transform 1 0 7084 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_46
timestamp 1618216021
transform 1 0 5336 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_50
timestamp 1618216021
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1618216021
transform 1 0 6716 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1618216021
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_69
timestamp 1618216021
transform 1 0 7452 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_81
timestamp 1618216021
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1618216021
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_87
timestamp 1618216021
transform 1 0 9108 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0803_
timestamp 1618216021
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0853_
timestamp 1618216021
transform 1 0 9752 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1618216021
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_101
timestamp 1618216021
transform 1 0 10396 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_105
timestamp 1618216021
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1618216021
transform 1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1618216021
transform 1 0 12972 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_i_clk
timestamp 1618216021
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_110
timestamp 1618216021
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1618216021
transform 1 0 11868 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1618216021
transform 1 0 12512 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1618216021
transform 1 0 12880 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1618216021
transform 1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1618216021
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1618216021
transform 1 0 13248 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_140
timestamp 1618216021
transform 1 0 13984 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1618216021
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_148
timestamp 1618216021
transform 1 0 14720 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1618216021
transform 1 0 15088 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0793_
timestamp 1618216021
transform 1 0 15456 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0794_
timestamp 1618216021
transform 1 0 16468 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1618216021
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1618216021
transform 1 0 17664 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1618216021
transform 1 0 18308 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1618216021
transform 1 0 17296 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1618216021
transform 1 0 17940 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_190
timestamp 1618216021
transform 1 0 18584 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1618216021
transform 1 0 20608 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1618216021
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1618216021
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_201
timestamp 1618216021
transform 1 0 19596 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_209
timestamp 1618216021
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1618216021
transform 1 0 22448 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0888_
timestamp 1618216021
transform 1 0 23092 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1618216021
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_235
timestamp 1618216021
transform 1 0 22724 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1618216021
transform 1 0 24104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0840_
timestamp 1618216021
transform 1 0 25208 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1618216021
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_246
timestamp 1618216021
transform 1 0 23736 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1618216021
transform 1 0 24380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1618216021
transform 1 0 24840 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1618216021
transform 1 0 26680 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_269
timestamp 1618216021
transform 1 0 25852 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_277
timestamp 1618216021
transform 1 0 26588 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_282
timestamp 1618216021
transform 1 0 27048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1618216021
transform -1 0 28428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1618216021
transform 1 0 27416 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1618216021
transform 1 0 27784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1618216021
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1618216021
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1618216021
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1618216021
transform 1 0 2024 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_6
timestamp 1618216021
transform 1 0 1656 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1618216021
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1618216021
transform 1 0 2300 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1618216021
transform 1 0 2944 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1618216021
transform 1 0 1472 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1618216021
transform 1 0 2852 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1618216021
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1618216021
transform 1 0 4232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1618216021
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1618216021
transform 1 0 4324 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_42
timestamp 1618216021
transform 1 0 4968 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1618216021
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_30
timestamp 1618216021
transform 1 0 3864 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_37
timestamp 1618216021
transform 1 0 4508 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_43
timestamp 1618216021
transform 1 0 5060 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0814_
timestamp 1618216021
transform 1 0 5336 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1618216021
transform 1 0 5152 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1178_
timestamp 1618216021
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1618216021
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_53
timestamp 1618216021
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_58
timestamp 1618216021
transform 1 0 6440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_60
timestamp 1618216021
transform 1 0 6624 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0596_
timestamp 1618216021
transform 1 0 7268 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1618216021
transform 1 0 7176 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1618216021
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1618216021
transform 1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_74
timestamp 1618216021
transform 1 0 7912 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_81
timestamp 1618216021
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1618216021
transform 1 0 8648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1618216021
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_85
timestamp 1618216021
transform 1 0 8924 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1618216021
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1618216021
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0534_
timestamp 1618216021
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0554_
timestamp 1618216021
transform 1 0 10672 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0848_
timestamp 1618216021
transform 1 0 9476 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0852_
timestamp 1618216021
transform 1 0 10212 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1618216021
transform 1 0 10304 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_108
timestamp 1618216021
transform 1 0 11040 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_95
timestamp 1618216021
transform 1 0 9844 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1618216021
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1618216021
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1618216021
transform 1 0 11224 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1618216021
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1618216021
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_122
timestamp 1618216021
transform 1 0 12328 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_126
timestamp 1618216021
transform 1 0 12696 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0546_
timestamp 1618216021
transform 1 0 13800 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1618216021
transform 1 0 14720 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1618216021
transform 1 0 14536 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1618216021
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1618216021
transform 1 0 13432 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1618216021
transform 1 0 14168 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_138
timestamp 1618216021
transform 1 0 13800 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1618216021
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1618216021
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0992_
timestamp 1618216021
transform 1 0 17112 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1618216021
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_162
timestamp 1618216021
transform 1 0 16008 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_170
timestamp 1618216021
transform 1 0 16744 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1618216021
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_164
timestamp 1618216021
transform 1 0 16192 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 1618216021
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0510_
timestamp 1618216021
transform 1 0 18308 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0516_
timestamp 1618216021
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1618216021
transform 1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _0795_
timestamp 1618216021
transform 1 0 17296 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_19_183
timestamp 1618216021
transform 1 0 17940 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_190
timestamp 1618216021
transform 1 0 18584 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1618216021
transform 1 0 17756 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_189
timestamp 1618216021
transform 1 0 18492 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_196
timestamp 1618216021
transform 1 0 19136 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0837_
timestamp 1618216021
transform 1 0 19964 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1618216021
transform 1 0 19504 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1618216021
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_198
timestamp 1618216021
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1618216021
transform 1 0 19872 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_201
timestamp 1618216021
transform 1 0 19596 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_209
timestamp 1618216021
transform 1 0 20332 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1618216021
transform 1 0 20884 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _0738_
timestamp 1618216021
transform 1 0 20976 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1618216021
transform 1 0 20240 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1618216021
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_224
timestamp 1618216021
transform 1 0 21712 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_229
timestamp 1618216021
transform 1 0 22172 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1618216021
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1618216021
transform 1 0 22448 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1618216021
transform 1 0 22908 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1618216021
transform 1 0 22724 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1618216021
transform 1 0 23092 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _0747_
timestamp 1618216021
transform 1 0 23184 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1618216021
transform 1 0 23000 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1618216021
transform 1 0 25116 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1618216021
transform 1 0 25208 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1618216021
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_254
timestamp 1618216021
transform 1 0 24472 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_260
timestamp 1618216021
transform 1 0 25024 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_252
timestamp 1618216021
transform 1 0 24288 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_256
timestamp 1618216021
transform 1 0 24656 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1618216021
transform 1 0 24840 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1031_
timestamp 1618216021
transform 1 0 27048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1618216021
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_278
timestamp 1618216021
transform 1 0 26680 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1618216021
transform -1 0 28428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1618216021
transform -1 0 28428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1618216021
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_286
timestamp 1618216021
transform 1 0 27416 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_286
timestamp 1618216021
transform 1 0 27416 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0960_
timestamp 1618216021
transform 1 0 1932 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1618216021
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1618216021
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_16
timestamp 1618216021
transform 1 0 2576 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0861_
timestamp 1618216021
transform 1 0 3496 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1618216021
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_33
timestamp 1618216021
transform 1 0 4140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0857_
timestamp 1618216021
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0862_
timestamp 1618216021
transform 1 0 5336 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1618216021
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_45
timestamp 1618216021
transform 1 0 5244 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1618216021
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_58
timestamp 1618216021
transform 1 0 6440 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1082_
timestamp 1618216021
transform 1 0 7544 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_21_66
timestamp 1618216021
transform 1 0 7176 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_87
timestamp 1618216021
transform 1 0 9108 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0851_
timestamp 1618216021
transform 1 0 9844 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0951_
timestamp 1618216021
transform 1 0 10580 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1618216021
transform 1 0 10212 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1089_
timestamp 1618216021
transform 1 0 12052 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1618216021
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_110
timestamp 1618216021
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1618216021
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0530_
timestamp 1618216021
transform 1 0 13984 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0845_
timestamp 1618216021
transform 1 0 14720 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1618216021
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1618216021
transform 1 0 14352 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0614_
timestamp 1618216021
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1618216021
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_155
timestamp 1618216021
transform 1 0 15364 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1618216021
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_172
timestamp 1618216021
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1059_
timestamp 1618216021
transform 1 0 17848 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_21_180
timestamp 1618216021
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o221ai_2  _0785_
timestamp 1618216021
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_199
timestamp 1618216021
transform 1 0 19412 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1618216021
transform 1 0 20884 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1618216021
transform 1 0 21252 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1618216021
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_223
timestamp 1618216021
transform 1 0 21620 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_227
timestamp 1618216021
transform 1 0 21988 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1618216021
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0757_
timestamp 1618216021
transform 1 0 24380 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1618216021
transform 1 0 23368 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_241
timestamp 1618216021
transform 1 0 23276 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1618216021
transform 1 0 24012 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_260
timestamp 1618216021
transform 1 0 25024 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1045_
timestamp 1618216021
transform 1 0 26588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1618216021
transform 1 0 25852 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_268
timestamp 1618216021
transform 1 0 25760 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_273
timestamp 1618216021
transform 1 0 26220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1618216021
transform 1 0 26956 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1618216021
transform -1 0 28428 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1618216021
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_286
timestamp 1618216021
transform 1 0 27416 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1618216021
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output157
timestamp 1618216021
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1618216021
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1618216021
transform 1 0 2116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _0533_
timestamp 1618216021
transform 1 0 4692 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1618216021
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_23
timestamp 1618216021
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_30
timestamp 1618216021
transform 1 0 3864 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_38
timestamp 1618216021
transform 1 0 4600 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0858_
timestamp 1618216021
transform 1 0 5796 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0961_
timestamp 1618216021
transform 1 0 6992 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_22_45
timestamp 1618216021
transform 1 0 5244 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_55
timestamp 1618216021
transform 1 0 6164 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_63
timestamp 1618216021
transform 1 0 6900 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0958_
timestamp 1618216021
transform 1 0 8004 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1618216021
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1618216021
transform 1 0 7636 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_82
timestamp 1618216021
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1618216021
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0952_
timestamp 1618216021
transform 1 0 10212 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1618216021
transform 1 0 9476 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1618216021
transform 1 0 9844 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1618216021
transform 1 0 10856 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1618216021
transform 1 0 11224 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_22_127
timestamp 1618216021
transform 1 0 12788 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1618216021
transform 1 0 13616 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0893_
timestamp 1618216021
transform 1 0 14720 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1618216021
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp 1618216021
transform 1 0 13524 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_139
timestamp 1618216021
transform 1 0 13892 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1618216021
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0784_
timestamp 1618216021
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0949_
timestamp 1618216021
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_155
timestamp 1618216021
transform 1 0 15364 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1618216021
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0706_
timestamp 1618216021
transform 1 0 18032 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1618216021
transform 1 0 17664 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_190
timestamp 1618216021
transform 1 0 18584 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0838_
timestamp 1618216021
transform 1 0 19964 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1618216021
transform 1 0 20976 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1618216021
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1618216021
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_201
timestamp 1618216021
transform 1 0 19596 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_209
timestamp 1618216021
transform 1 0 20332 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_215
timestamp 1618216021
transform 1 0 20884 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_232
timestamp 1618216021
transform 1 0 22448 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1618216021
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_244
timestamp 1618216021
transform 1 0 23552 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_256
timestamp 1618216021
transform 1 0 24656 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1618216021
transform 1 0 24840 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_262
timestamp 1618216021
transform 1 0 25208 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0624_
timestamp 1618216021
transform 1 0 25300 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1618216021
transform 1 0 26312 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1618216021
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1618216021
transform -1 0 28428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_290
timestamp 1618216021
transform 1 0 27784 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1618216021
transform 1 0 2944 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1618216021
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1618216021
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_6
timestamp 1618216021
transform 1 0 1656 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_18
timestamp 1618216021
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1618216021
transform 1 0 4416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1618216021
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1618216021
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_48
timestamp 1618216021
transform 1 0 5520 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_56
timestamp 1618216021
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1618216021
transform 1 0 6440 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1618216021
transform 1 0 7084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_4  _0597_
timestamp 1618216021
transform 1 0 8096 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_23_73
timestamp 1618216021
transform 1 0 7820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0581_
timestamp 1618216021
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1618216021
transform 1 0 10028 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_105
timestamp 1618216021
transform 1 0 10764 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0947_
timestamp 1618216021
transform 1 0 12052 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1618216021
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1618216021
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1618216021
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1618216021
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1618216021
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0847_
timestamp 1618216021
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0892_
timestamp 1618216021
transform 1 0 14720 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_23_134
timestamp 1618216021
transform 1 0 13432 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1618216021
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0850_
timestamp 1618216021
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1618216021
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1618216021
transform 1 0 15364 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1618216021
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1618216021
transform 1 0 16928 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1618216021
transform 1 0 18492 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0783_
timestamp 1618216021
transform 1 0 17296 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_23_183
timestamp 1618216021
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_192
timestamp 1618216021
transform 1 0 18768 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp 1618216021
transform 1 0 21068 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0776_
timestamp 1618216021
transform 1 0 19688 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1618216021
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_209
timestamp 1618216021
transform 1 0 20332 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0765_
timestamp 1618216021
transform 1 0 22816 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1618216021
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_224
timestamp 1618216021
transform 1 0 21712 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_229
timestamp 1618216021
transform 1 0 22172 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_235
timestamp 1618216021
transform 1 0 22724 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0748_
timestamp 1618216021
transform 1 0 23920 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1618216021
transform 1 0 23460 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1618216021
transform 1 0 23828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_255
timestamp 1618216021
transform 1 0 24564 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp 1618216021
transform 1 0 25484 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_263
timestamp 1618216021
transform 1 0 25300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1618216021
transform 1 0 26956 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1618216021
transform -1 0 28428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1618216021
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_286
timestamp 1618216021
transform 1 0 27416 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1618216021
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1618216021
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_6
timestamp 1618216021
transform 1 0 1656 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1618216021
transform 1 0 2760 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1618216021
transform 1 0 4232 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1618216021
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_26
timestamp 1618216021
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_30
timestamp 1618216021
transform 1 0 3864 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0864_
timestamp 1618216021
transform 1 0 6532 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_50
timestamp 1618216021
transform 1 0 5704 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_58
timestamp 1618216021
transform 1 0 6440 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_63
timestamp 1618216021
transform 1 0 6900 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0896_
timestamp 1618216021
transform 1 0 7268 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0957_
timestamp 1618216021
transform 1 0 8280 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1618216021
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_71
timestamp 1618216021
transform 1 0 7636 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_77
timestamp 1618216021
transform 1 0 8188 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_82
timestamp 1618216021
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1618216021
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0589_
timestamp 1618216021
transform 1 0 9476 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0950_
timestamp 1618216021
transform 1 0 10764 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_98
timestamp 1618216021
transform 1 0 10120 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_104
timestamp 1618216021
transform 1 0 10672 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1618216021
transform 1 0 11132 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _1012_
timestamp 1618216021
transform 1 0 13156 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1618216021
transform 1 0 12236 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1618216021
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1618216021
transform 1 0 14720 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1618216021
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_138
timestamp 1618216021
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1618216021
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1618216021
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0946_
timestamp 1618216021
transform 1 0 16744 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_164
timestamp 1618216021
transform 1 0 16192 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_174
timestamp 1618216021
transform 1 0 17112 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1618216021
transform 1 0 17480 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1618216021
transform 1 0 18124 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1618216021
transform 1 0 18768 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1618216021
transform 1 0 17756 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_188
timestamp 1618216021
transform 1 0 18400 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_195
timestamp 1618216021
transform 1 0 19044 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1618216021
transform 1 0 19964 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1618216021
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1618216021
transform 1 0 19412 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1618216021
transform 1 0 19596 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0740_
timestamp 1618216021
transform 1 0 21804 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1190_
timestamp 1618216021
transform 1 0 22540 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1618216021
transform 1 0 21436 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_229
timestamp 1618216021
transform 1 0 22172 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1618216021
transform 1 0 25208 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1618216021
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_250
timestamp 1618216021
transform 1 0 24104 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_256
timestamp 1618216021
transform 1 0 24656 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1618216021
transform 1 0 24840 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0598_
timestamp 1618216021
transform 1 0 27048 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_278
timestamp 1618216021
transform 1 0 26680 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1618216021
transform -1 0 28428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp 1618216021
transform 1 0 27692 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_293
timestamp 1618216021
transform 1 0 28060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1039_
timestamp 1618216021
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1618216021
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1618216021
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1618216021
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0901_
timestamp 1618216021
transform 1 0 3588 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0904_
timestamp 1618216021
transform 1 0 4600 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1618216021
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0865_
timestamp 1618216021
transform 1 0 5612 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0869_
timestamp 1618216021
transform 1 0 6808 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1618216021
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 1618216021
transform 1 0 5244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1618216021
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1618216021
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1618216021
transform 1 0 8464 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1618216021
transform 1 0 7452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_77
timestamp 1618216021
transform 1 0 8188 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_97
timestamp 1618216021
transform 1 0 10028 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1618216021
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1618216021
transform 1 0 12052 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1618216021
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1618216021
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1618216021
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1618216021
transform 1 0 13892 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_clk
timestamp 1618216021
transform 1 0 14628 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1618216021
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1618216021
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_146
timestamp 1618216021
transform 1 0 14536 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1618216021
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_167
timestamp 1618216021
transform 1 0 16468 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1618216021
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1618216021
transform 1 0 18860 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0991_
timestamp 1618216021
transform 1 0 17296 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_25_183
timestamp 1618216021
transform 1 0 17940 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1618216021
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1618216021
transform 1 0 19136 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1618216021
transform 1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_203
timestamp 1618216021
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1618216021
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0654_
timestamp 1618216021
transform 1 0 22540 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0695_
timestamp 1618216021
transform 1 0 21344 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1618216021
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1618216021
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_224
timestamp 1618216021
transform 1 0 21712 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_229
timestamp 1618216021
transform 1 0 22172 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1618216021
transform 1 0 22908 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0749_
timestamp 1618216021
transform 1 0 23276 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1618216021
transform 1 0 24564 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1618216021
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_253
timestamp 1618216021
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1618216021
transform 1 0 26588 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_271
timestamp 1618216021
transform 1 0 26036 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1618216021
transform 1 0 26956 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1618216021
transform -1 0 28428 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1618216021
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_286
timestamp 1618216021
transform 1 0 27416 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0968_
timestamp 1618216021
transform 1 0 2484 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1077_
timestamp 1618216021
transform 1 0 1656 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1618216021
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1618216021
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1618216021
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_6
timestamp 1618216021
transform 1 0 1656 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_14
timestamp 1618216021
transform 1 0 2392 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1618216021
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0969_
timestamp 1618216021
transform 1 0 3588 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1618216021
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1618216021
transform 1 0 3128 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1618216021
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_30
timestamp 1618216021
transform 1 0 3864 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1618216021
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1618216021
transform 1 0 4600 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1618216021
transform 1 0 4232 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1618216021
transform 1 0 4232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_41
timestamp 1618216021
transform 1 0 4876 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_37
timestamp 1618216021
transform 1 0 4508 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o211ai_2  _0638_
timestamp 1618216021
transform 1 0 7084 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0817_
timestamp 1618216021
transform 1 0 5612 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1618216021
transform 1 0 5888 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1618216021
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_49
timestamp 1618216021
transform 1 0 5612 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_53
timestamp 1618216021
transform 1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_58
timestamp 1618216021
transform 1 0 6440 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_64
timestamp 1618216021
transform 1 0 6992 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1618216021
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1618216021
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1618216021
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1618216021
transform 1 0 7360 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1618216021
transform 1 0 8004 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_83
timestamp 1618216021
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1618216021
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_75
timestamp 1618216021
transform 1 0 8004 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1618216021
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _0963_
timestamp 1618216021
transform 1 0 9660 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp 1618216021
transform 1 0 9476 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1618216021
transform 1 0 10948 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_89
timestamp 1618216021
transform 1 0 9292 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_97
timestamp 1618216021
transform 1 0 10028 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_109
timestamp 1618216021
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0625_
timestamp 1618216021
transform 1 0 11316 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1618216021
transform 1 0 12420 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1618216021
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_115
timestamp 1618216021
transform 1 0 11684 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_130
timestamp 1618216021
transform 1 0 13064 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1618216021
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1618216021
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_127
timestamp 1618216021
transform 1 0 12788 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0508_
timestamp 1618216021
transform 1 0 14260 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0540_
timestamp 1618216021
transform 1 0 13524 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1618216021
transform 1 0 14720 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1618216021
transform 1 0 14996 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1618216021
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1618216021
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1618216021
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1618216021
transform 1 0 13892 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1618216021
transform 1 0 14628 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1618216021
transform 1 0 15732 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1618216021
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1618216021
transform 1 0 15364 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_167
timestamp 1618216021
transform 1 0 16468 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1618216021
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1618216021
transform 1 0 17296 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1060_
timestamp 1618216021
transform 1 0 17572 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1618216021
transform 1 0 17204 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1618216021
transform 1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_185
timestamp 1618216021
transform 1 0 18124 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0712_
timestamp 1618216021
transform 1 0 20332 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1618216021
transform 1 0 20148 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1618216021
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_201
timestamp 1618216021
transform 1 0 19596 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_197
timestamp 1618216021
transform 1 0 19228 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_216
timestamp 1618216021
transform 1 0 20976 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0639_
timestamp 1618216021
transform 1 0 22540 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1618216021
transform 1 0 22540 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1618216021
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_223
timestamp 1618216021
transform 1 0 21620 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1618216021
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_229
timestamp 1618216021
transform 1 0 22172 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_240
timestamp 1618216021
transform 1 0 23184 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0632_
timestamp 1618216021
transform 1 0 25024 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1618216021
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_249
timestamp 1618216021
transform 1 0 24012 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1618216021
transform 1 0 24840 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_252
timestamp 1618216021
transform 1 0 24288 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1043_
timestamp 1618216021
transform 1 0 26956 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1618216021
transform 1 0 25576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1618216021
transform 1 0 26588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1618216021
transform 1 0 26220 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_269
timestamp 1618216021
transform 1 0 25852 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1618216021
transform 1 0 26588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_267
timestamp 1618216021
transform 1 0 25668 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1618216021
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1618216021
transform 1 0 26956 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1618216021
transform -1 0 28428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1618216021
transform -1 0 28428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1618216021
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_285
timestamp 1618216021
transform 1 0 27324 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_293
timestamp 1618216021
transform 1 0 28060 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_286
timestamp 1618216021
transform 1 0 27416 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1618216021
transform 1 0 1564 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1618216021
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1618216021
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_21
timestamp 1618216021
transform 1 0 3036 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0822_
timestamp 1618216021
transform 1 0 4232 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1618216021
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_30
timestamp 1618216021
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1618216021
transform 1 0 4876 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1618216021
transform 1 0 5704 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_49
timestamp 1618216021
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1618216021
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0816_
timestamp 1618216021
transform 1 0 7544 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1618216021
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1618216021
transform 1 0 7176 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1618216021
transform 1 0 7912 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_81
timestamp 1618216021
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1618216021
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_87
timestamp 1618216021
transform 1 0 9108 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0646_
timestamp 1618216021
transform 1 0 9936 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_28_95
timestamp 1618216021
transform 1 0 9844 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_103
timestamp 1618216021
transform 1 0 10580 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1618216021
transform 1 0 11500 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1618216021
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_129
timestamp 1618216021
transform 1 0 12972 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0525_
timestamp 1618216021
transform 1 0 13616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0677_
timestamp 1618216021
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1618216021
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_135
timestamp 1618216021
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1618216021
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1618216021
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1618216021
transform 1 0 15088 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0799_
timestamp 1618216021
transform 1 0 15456 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0802_
timestamp 1618216021
transform 1 0 16192 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1618216021
transform 1 0 15824 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1618216021
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_i_clk
timestamp 1618216021
transform 1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1618216021
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_192
timestamp 1618216021
transform 1 0 18768 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_196
timestamp 1618216021
transform 1 0 19136 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1618216021
transform 1 0 19964 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1618216021
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_201
timestamp 1618216021
transform 1 0 19596 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_208
timestamp 1618216021
transform 1 0 20240 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0704_
timestamp 1618216021
transform 1 0 21988 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_220
timestamp 1618216021
transform 1 0 21344 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_226
timestamp 1618216021
transform 1 0 21896 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_231
timestamp 1618216021
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1618216021
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1618216021
transform 1 0 25208 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_243
timestamp 1618216021
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_255
timestamp 1618216021
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1618216021
transform 1 0 24840 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1618216021
transform 1 0 25944 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_266
timestamp 1618216021
transform 1 0 25576 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1618216021
transform -1 0 28428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_286
timestamp 1618216021
transform 1 0 27416 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1040_
timestamp 1618216021
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1618216021
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1618216021
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1618216021
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp 1618216021
transform 1 0 2484 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_21
timestamp 1618216021
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1618216021
transform 1 0 3128 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_38
timestamp 1618216021
transform 1 0 4600 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _0623_
timestamp 1618216021
transform 1 0 6808 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0870_
timestamp 1618216021
transform 1 0 5336 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1618216021
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_53
timestamp 1618216021
transform 1 0 5980 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_58
timestamp 1618216021
transform 1 0 6440 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_79
timestamp 1618216021
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp 1618216021
transform 1 0 9568 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_91
timestamp 1618216021
transform 1 0 9476 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_108
timestamp 1618216021
transform 1 0 11040 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1618216021
transform 1 0 13064 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0653_
timestamp 1618216021
transform 1 0 12052 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1618216021
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1618216021
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1618216021
transform 1 0 12696 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0507_
timestamp 1618216021
transform 1 0 13892 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _0770_
timestamp 1618216021
transform 1 0 14628 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_133
timestamp 1618216021
transform 1 0 13340 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_143
timestamp 1618216021
transform 1 0 14260 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1618216021
transform 1 0 15824 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1618216021
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_156
timestamp 1618216021
transform 1 0 15456 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_164
timestamp 1618216021
transform 1 0 16192 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_170
timestamp 1618216021
transform 1 0 16744 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1618216021
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0574_
timestamp 1618216021
transform 1 0 17756 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0697_
timestamp 1618216021
transform 1 0 18676 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_180
timestamp 1618216021
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_187
timestamp 1618216021
transform 1 0 18308 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0824_
timestamp 1618216021
transform 1 0 20976 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0825_
timestamp 1618216021
transform 1 0 19964 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_29_197
timestamp 1618216021
transform 1 0 19228 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_212
timestamp 1618216021
transform 1 0 20608 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1618216021
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_i_clk
timestamp 1618216021
transform 1 0 22632 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_219
timestamp 1618216021
transform 1 0 21252 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_227
timestamp 1618216021
transform 1 0 21988 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1618216021
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 1618216021
transform 1 0 22540 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_237
timestamp 1618216021
transform 1 0 22908 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_i_clk
timestamp 1618216021
transform 1 0 23736 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_245
timestamp 1618216021
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1618216021
transform 1 0 24012 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_261
timestamp 1618216021
transform 1 0 25116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1618216021
transform 1 0 25392 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_280
timestamp 1618216021
transform 1 0 26864 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1618216021
transform -1 0 28428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1618216021
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_284
timestamp 1618216021
transform 1 0 27232 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_286
timestamp 1618216021
transform 1 0 27416 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1046_
timestamp 1618216021
transform 1 0 2116 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1618216021
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1618216021
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_7
timestamp 1618216021
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1618216021
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0821_
timestamp 1618216021
transform 1 0 4232 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1618216021
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1618216021
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_30
timestamp 1618216021
transform 1 0 3864 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1618216021
transform 1 0 4876 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1618216021
transform 1 0 5244 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0637_
timestamp 1618216021
transform 1 0 5980 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_48
timestamp 1618216021
transform 1 0 5520 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_52
timestamp 1618216021
transform 1 0 5888 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1618216021
transform 1 0 6808 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _0645_
timestamp 1618216021
transform 1 0 8004 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1618216021
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_i_clk
timestamp 1618216021
transform 1 0 7176 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_69
timestamp 1618216021
transform 1 0 7452 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_81
timestamp 1618216021
transform 1 0 8556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1618216021
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1618216021
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0522_
timestamp 1618216021
transform 1 0 9476 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0592_
timestamp 1618216021
transform 1 0 10396 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1618216021
transform 1 0 10028 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_107
timestamp 1618216021
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0520_
timestamp 1618216021
transform 1 0 12972 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0527_
timestamp 1618216021
transform 1 0 11776 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1618216021
transform 1 0 11684 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_120
timestamp 1618216021
transform 1 0 12144 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_128
timestamp 1618216021
transform 1 0 12880 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0726_
timestamp 1618216021
transform 1 0 14720 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1618216021
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_134
timestamp 1618216021
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1618216021
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1618216021
transform 1 0 14352 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1618216021
transform 1 0 17112 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0993_
timestamp 1618216021
transform 1 0 15916 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1618216021
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1618216021
transform 1 0 16744 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0652_
timestamp 1618216021
transform 1 0 17756 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1618216021
transform 1 0 17388 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_193
timestamp 1618216021
transform 1 0 18860 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1618216021
transform 1 0 19964 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1618216021
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1618216021
transform 1 0 19412 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1618216021
transform 1 0 19596 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1618216021
transform 1 0 22724 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1618216021
transform 1 0 21436 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_233
timestamp 1618216021
transform 1 0 22540 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1618216021
transform 1 0 24104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0662_
timestamp 1618216021
transform 1 0 25208 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1618216021
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1618216021
transform 1 0 23368 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1618216021
transform 1 0 24380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1618216021
transform 1 0 24840 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0672_
timestamp 1618216021
transform 1 0 26220 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_269
timestamp 1618216021
transform 1 0 25852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_280
timestamp 1618216021
transform 1 0 26864 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1618216021
transform -1 0 28428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1618216021
transform 1 0 27416 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1618216021
transform 1 0 27784 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1618216021
transform 1 0 3036 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1618216021
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1618216021
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_15
timestamp 1618216021
transform 1 0 2484 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1618216021
transform 1 0 5060 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_37
timestamp 1618216021
transform 1 0 4508 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1618216021
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0644_
timestamp 1618216021
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1618216021
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_46
timestamp 1618216021
transform 1 0 5336 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_53
timestamp 1618216021
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_58
timestamp 1618216021
transform 1 0 6440 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1618216021
transform 1 0 8740 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_71
timestamp 1618216021
transform 1 0 7636 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_86
timestamp 1618216021
transform 1 0 9016 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0532_
timestamp 1618216021
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1618216021
transform 1 0 9568 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_i_clk
timestamp 1618216021
transform 1 0 10948 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp 1618216021
transform 1 0 9844 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1618216021
transform 1 0 10580 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0666_
timestamp 1618216021
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1618216021
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_110
timestamp 1618216021
transform 1 0 11224 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_115
timestamp 1618216021
transform 1 0 11684 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_129
timestamp 1618216021
transform 1 0 12972 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0515_
timestamp 1618216021
transform 1 0 13708 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0521_
timestamp 1618216021
transform 1 0 14904 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1618216021
transform 1 0 14536 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1618216021
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1618216021
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1618216021
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1618216021
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_166
timestamp 1618216021
transform 1 0 16376 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_170
timestamp 1618216021
transform 1 0 16744 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1618216021
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1618216021
transform 1 0 17296 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1618216021
transform 1 0 19044 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_185
timestamp 1618216021
transform 1 0 18124 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1618216021
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _0826_
timestamp 1618216021
transform 1 0 20884 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1618216021
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1618216021
transform 1 0 22908 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1618216021
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_222
timestamp 1618216021
transform 1 0 21528 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_229
timestamp 1618216021
transform 1 0 22172 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1618216021
transform 1 0 24748 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_253
timestamp 1618216021
transform 1 0 24380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1028_
timestamp 1618216021
transform 1 0 26588 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_273
timestamp 1618216021
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1618216021
transform 1 0 26956 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1618216021
transform -1 0 28428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1618216021
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_286
timestamp 1618216021
transform 1 0 27416 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0966_
timestamp 1618216021
transform 1 0 2392 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1618216021
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1618216021
transform 1 0 1656 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1618216021
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_10
timestamp 1618216021
transform 1 0 2024 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_21
timestamp 1618216021
transform 1 0 3036 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1618216021
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1618216021
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_42
timestamp 1618216021
transform 1 0 4968 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0818_
timestamp 1618216021
transform 1 0 6900 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0867_
timestamp 1618216021
transform 1 0 5244 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_i_clk
timestamp 1618216021
transform 1 0 6256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_52
timestamp 1618216021
transform 1 0 5888 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_59
timestamp 1618216021
transform 1 0 6532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1618216021
transform 1 0 8188 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1618216021
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_70
timestamp 1618216021
transform 1 0 7544 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_76
timestamp 1618216021
transform 1 0 8096 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_80
timestamp 1618216021
transform 1 0 8464 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_87
timestamp 1618216021
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_4  _0612_
timestamp 1618216021
transform 1 0 9476 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__or4_4  _0531_
timestamp 1618216021
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0617_
timestamp 1618216021
transform 1 0 11776 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1618216021
transform 1 0 11408 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_120
timestamp 1618216021
transform 1 0 12144 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1618216021
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0526_
timestamp 1618216021
transform 1 0 14720 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1618216021
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_139
timestamp 1618216021
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1618216021
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1056_
timestamp 1618216021
transform 1 0 16192 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_32_157
timestamp 1618216021
transform 1 0 15548 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_163
timestamp 1618216021
transform 1 0 16100 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0656_
timestamp 1618216021
transform 1 0 18124 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1618216021
transform 1 0 17756 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_191
timestamp 1618216021
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0823_
timestamp 1618216021
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1618216021
transform 1 0 20700 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1618216021
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1618216021
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1618216021
transform 1 0 19596 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1618216021
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0827_
timestamp 1618216021
transform 1 0 22816 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_32_229
timestamp 1618216021
transform 1 0 22172 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_235
timestamp 1618216021
transform 1 0 22724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0663_
timestamp 1618216021
transform 1 0 23828 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1618216021
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_243
timestamp 1618216021
transform 1 0 23460 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_251
timestamp 1618216021
transform 1 0 24196 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_258
timestamp 1618216021
transform 1 0 24840 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 1618216021
transform 1 0 25760 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_266
timestamp 1618216021
transform 1 0 25576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1618216021
transform -1 0 28428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_284
timestamp 1618216021
transform 1 0 27232 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_292
timestamp 1618216021
transform 1 0 27968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _0819_
timestamp 1618216021
transform 1 0 2760 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1079_
timestamp 1618216021
transform 1 0 1564 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1618216021
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1618216021
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output151
timestamp 1618216021
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1618216021
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1618216021
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_11
timestamp 1618216021
transform 1 0 2116 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_17
timestamp 1618216021
transform 1 0 2668 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1618216021
transform 1 0 3496 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1618216021
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1618216021
transform 1 0 3128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_29
timestamp 1618216021
transform 1 0 3772 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_25
timestamp 1618216021
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_30
timestamp 1618216021
transform 1 0 3864 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0622_
timestamp 1618216021
transform 1 0 4692 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1618216021
transform 1 0 4140 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_38
timestamp 1618216021
transform 1 0 4600 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1618216021
transform 1 0 4232 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1618216021
transform 1 0 5888 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1618216021
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1618216021
transform 1 0 5704 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_56
timestamp 1618216021
transform 1 0 6256 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_58
timestamp 1618216021
transform 1 0 6440 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_48
timestamp 1618216021
transform 1 0 5520 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0611_
timestamp 1618216021
transform 1 0 8004 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1618216021
transform 1 0 7176 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1618216021
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_82
timestamp 1618216021
transform 1 0 8648 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_68
timestamp 1618216021
transform 1 0 7360 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_74
timestamp 1618216021
transform 1 0 7912 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_82
timestamp 1618216021
transform 1 0 8648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1618216021
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1618216021
transform 1 0 9476 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0631_
timestamp 1618216021
transform 1 0 9292 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _1078_
timestamp 1618216021
transform 1 0 10396 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_33_88
timestamp 1618216021
transform 1 0 9200 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_94
timestamp 1618216021
transform 1 0 9752 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_100
timestamp 1618216021
transform 1 0 10304 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1618216021
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_110
timestamp 1618216021
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_115
timestamp 1618216021
transform 1 0 11684 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1618216021
transform 1 0 11960 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0610_
timestamp 1618216021
transform 1 0 12236 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0619_
timestamp 1618216021
transform 1 0 12328 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1618216021
transform 1 0 12604 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_126
timestamp 1618216021
transform 1 0 12696 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0543_
timestamp 1618216021
transform 1 0 12972 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0944_
timestamp 1618216021
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0529_
timestamp 1618216021
transform 1 0 13708 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0798_
timestamp 1618216021
transform 1 0 14720 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _1007_
timestamp 1618216021
transform 1 0 14996 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1618216021
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1618216021
transform 1 0 13340 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1618216021
transform 1 0 14536 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1618216021
transform 1 0 14904 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_139
timestamp 1618216021
transform 1 0 13892 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1618216021
transform 1 0 14352 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0668_
timestamp 1618216021
transform 1 0 15916 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0970_
timestamp 1618216021
transform 1 0 17112 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1618216021
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_164
timestamp 1618216021
transform 1 0 16192 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_170
timestamp 1618216021
transform 1 0 16744 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_172
timestamp 1618216021
transform 1 0 16928 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_157
timestamp 1618216021
transform 1 0 15548 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 1618216021
transform 1 0 16284 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_173
timestamp 1618216021
transform 1 0 17020 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0594_
timestamp 1618216021
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0651_
timestamp 1618216021
transform 1 0 17940 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _0661_
timestamp 1618216021
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1618216021
transform 1 0 17664 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1618216021
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1618216021
transform 1 0 17480 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_182
timestamp 1618216021
transform 1 0 17848 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_190
timestamp 1618216021
transform 1 0 18584 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1618216021
transform 1 0 19504 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0872_
timestamp 1618216021
transform 1 0 19964 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1618216021
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_203
timestamp 1618216021
transform 1 0 19780 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_198
timestamp 1618216021
transform 1 0 19320 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1618216021
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1618216021
transform 1 0 20700 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0829_
timestamp 1618216021
transform 1 0 20608 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_33_211
timestamp 1618216021
transform 1 0 20516 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1618216021
transform 1 0 20332 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_216
timestamp 1618216021
transform 1 0 20976 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1618216021
transform 1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1618216021
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_219
timestamp 1618216021
transform 1 0 21252 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_227
timestamp 1618216021
transform 1 0 21988 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_229
timestamp 1618216021
transform 1 0 22172 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp 1618216021
transform 1 0 21712 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1618216021
transform 1 0 22080 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1618216021
transform 1 0 23184 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1618216021
transform 1 0 22540 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1618216021
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_232
timestamp 1618216021
transform 1 0 22448 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_236
timestamp 1618216021
transform 1 0 22816 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0671_
timestamp 1618216021
transform 1 0 23092 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1618216021
transform 1 0 23828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_243
timestamp 1618216021
transform 1 0 23460 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_251
timestamp 1618216021
transform 1 0 24196 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_250
timestamp 1618216021
transform 1 0 24104 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1618216021
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1618216021
transform 1 0 24748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_256
timestamp 1618216021
transform 1 0 24656 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1618216021
transform 1 0 24840 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp 1618216021
transform 1 0 25116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_262
timestamp 1618216021
transform 1 0 25208 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0975_
timestamp 1618216021
transform 1 0 25300 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1618216021
transform 1 0 26312 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1618216021
transform 1 0 25484 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1618216021
transform 1 0 26956 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1618216021
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1618216021
transform -1 0 28428 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1618216021
transform -1 0 28428 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1618216021
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_286
timestamp 1618216021
transform 1 0 27416 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1618216021
transform 1 0 27784 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1618216021
transform 1 0 2116 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1618216021
transform 1 0 2760 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1618216021
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1618216021
transform 1 0 1472 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1618216021
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1618216021
transform 1 0 1748 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1618216021
transform 1 0 2392 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1618216021
transform 1 0 4692 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1618216021
transform 1 0 4232 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_38
timestamp 1618216021
transform 1 0 4600 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_42
timestamp 1618216021
transform 1 0 4968 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0820_
timestamp 1618216021
transform 1 0 5336 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1618216021
transform 1 0 6808 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1618216021
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_53
timestamp 1618216021
transform 1 0 5980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_58
timestamp 1618216021
transform 1 0 6440 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0630_
timestamp 1618216021
transform 1 0 8648 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_78
timestamp 1618216021
transform 1 0 8280 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1618216021
transform 1 0 9660 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_89
timestamp 1618216021
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_109
timestamp 1618216021
transform 1 0 11132 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0519_
timestamp 1618216021
transform 1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0971_
timestamp 1618216021
transform 1 0 13156 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1618216021
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1618216021
transform 1 0 11500 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_115
timestamp 1618216021
transform 1 0 11684 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_123
timestamp 1618216021
transform 1 0 12420 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1618216021
transform 1 0 12788 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0846_
timestamp 1618216021
transform 1 0 13892 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0945_
timestamp 1618216021
transform 1 0 15088 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_135
timestamp 1618216021
transform 1 0 13524 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_148
timestamp 1618216021
transform 1 0 14720 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1618216021
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_161
timestamp 1618216021
transform 1 0 15916 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1618216021
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_172
timestamp 1618216021
transform 1 0 16928 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1618216021
transform 1 0 18860 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0660_
timestamp 1618216021
transform 1 0 17848 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_35_180
timestamp 1618216021
transform 1 0 17664 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1618216021
transform 1 0 18492 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1618216021
transform 1 0 19136 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1618216021
transform 1 0 19504 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_216
timestamp 1618216021
transform 1 0 20976 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1618216021
transform 1 0 21344 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0670_
timestamp 1618216021
transform 1 0 22540 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1618216021
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_223
timestamp 1618216021
transform 1 0 21620 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_227
timestamp 1618216021
transform 1 0 21988 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_229
timestamp 1618216021
transform 1 0 22172 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1618216021
transform 1 0 23184 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1618216021
transform 1 0 24656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0680_
timestamp 1618216021
transform 1 0 23644 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_35_244
timestamp 1618216021
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_252
timestamp 1618216021
transform 1 0 24288 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_259
timestamp 1618216021
transform 1 0 24932 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1618216021
transform 1 0 25300 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0972_
timestamp 1618216021
transform 1 0 25944 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_266
timestamp 1618216021
transform 1 0 25576 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1618216021
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1618216021
transform -1 0 28428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1618216021
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_286
timestamp 1618216021
transform 1 0 27416 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1618216021
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1618216021
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1618216021
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1618216021
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1618216021
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1618216021
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_42
timestamp 1618216021
transform 1 0 4968 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1618216021
transform 1 0 5612 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_36_48
timestamp 1618216021
transform 1 0 5520 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1618216021
transform 1 0 7084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1618216021
transform 1 0 7452 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1618216021
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1618216021
transform 1 0 8096 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1618216021
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1618216021
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1618216021
transform 1 0 10488 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0965_
timestamp 1618216021
transform 1 0 9476 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1618216021
transform 1 0 10120 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_105
timestamp 1618216021
transform 1 0 10764 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0834_
timestamp 1618216021
transform 1 0 11408 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_i_clk
timestamp 1618216021
transform 1 0 12420 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_111
timestamp 1618216021
transform 1 0 11316 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1618216021
transform 1 0 12052 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_126
timestamp 1618216021
transform 1 0 12696 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1618216021
transform 1 0 13432 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1618216021
transform 1 0 14720 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1618216021
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_137
timestamp 1618216021
transform 1 0 13708 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_144
timestamp 1618216021
transform 1 0 14352 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_151
timestamp 1618216021
transform 1 0 14996 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0830_
timestamp 1618216021
transform 1 0 15364 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1074_
timestamp 1618216021
transform 1 0 16192 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1618216021
transform 1 0 15732 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_163
timestamp 1618216021
transform 1 0 16100 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0874_
timestamp 1618216021
transform 1 0 18492 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_36_181
timestamp 1618216021
transform 1 0 17756 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_196
timestamp 1618216021
transform 1 0 19136 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0871_
timestamp 1618216021
transform 1 0 20976 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1618216021
transform 1 0 19964 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1618216021
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1618216021
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1618216021
transform 1 0 20608 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1618216021
transform 1 0 21804 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1618216021
transform 1 0 21344 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_224
timestamp 1618216021
transform 1 0 21712 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _0679_
timestamp 1618216021
transform 1 0 23644 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0974_
timestamp 1618216021
transform 1 0 25208 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1618216021
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_241
timestamp 1618216021
transform 1 0 23276 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_252
timestamp 1618216021
transform 1 0 24288 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_256
timestamp 1618216021
transform 1 0 24656 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_258
timestamp 1618216021
transform 1 0 24840 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output155
timestamp 1618216021
transform 1 0 26680 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_269
timestamp 1618216021
transform 1 0 25852 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_277
timestamp 1618216021
transform 1 0 26588 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_282
timestamp 1618216021
transform 1 0 27048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1618216021
transform -1 0 28428 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1618216021
transform 1 0 27416 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_290
timestamp 1618216021
transform 1 0 27784 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1618216021
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output133
timestamp 1618216021
transform 1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1618216021
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_11
timestamp 1618216021
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_23
timestamp 1618216021
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_35
timestamp 1618216021
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0866_
timestamp 1618216021
transform 1 0 6808 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1618216021
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_i_clk
timestamp 1618216021
transform 1 0 5704 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_47
timestamp 1618216021
transform 1 0 5428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_53
timestamp 1618216021
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_58
timestamp 1618216021
transform 1 0 6440 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1618216021
transform 1 0 8924 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1618216021
transform 1 0 7820 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_69
timestamp 1618216021
transform 1 0 7452 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_76
timestamp 1618216021
transform 1 0 8096 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_84
timestamp 1618216021
transform 1 0 8832 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0967_
timestamp 1618216021
transform 1 0 9844 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_i_clk
timestamp 1618216021
transform 1 0 10856 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_88
timestamp 1618216021
transform 1 0 9200 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_94
timestamp 1618216021
transform 1 0 9752 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_102
timestamp 1618216021
transform 1 0 10488 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_109
timestamp 1618216021
transform 1 0 11132 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1618216021
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1618216021
transform 1 0 12788 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1618216021
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1618216021
transform 1 0 11500 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_115
timestamp 1618216021
transform 1 0 11684 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_122
timestamp 1618216021
transform 1 0 12328 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_126
timestamp 1618216021
transform 1 0 12696 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0725_
timestamp 1618216021
transform 1 0 14628 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1618216021
transform 1 0 14260 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_151
timestamp 1618216021
transform 1 0 14996 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0831_
timestamp 1618216021
transform 1 0 16100 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0878_
timestamp 1618216021
transform 1 0 15364 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1618216021
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_159
timestamp 1618216021
transform 1 0 15732 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_167
timestamp 1618216021
transform 1 0 16468 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_172
timestamp 1618216021
transform 1 0 16928 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0973_
timestamp 1618216021
transform 1 0 17296 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1618216021
transform 1 0 18676 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_37_183
timestamp 1618216021
transform 1 0 17940 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0876_
timestamp 1618216021
transform 1 0 21068 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_37_207
timestamp 1618216021
transform 1 0 20148 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_215
timestamp 1618216021
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _0875_
timestamp 1618216021
transform 1 0 22540 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1618216021
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_224
timestamp 1618216021
transform 1 0 21712 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_229
timestamp 1618216021
transform 1 0 22172 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_240
timestamp 1618216021
transform 1 0 23184 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1073_
timestamp 1618216021
transform 1 0 24012 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_37_248
timestamp 1618216021
transform 1 0 23920 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1618216021
transform 1 0 25944 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1618216021
transform 1 0 26588 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1618216021
transform 1 0 25576 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_273
timestamp 1618216021
transform 1 0 26220 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1618216021
transform 1 0 26956 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1618216021
transform -1 0 28428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1618216021
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_286
timestamp 1618216021
transform 1 0 27416 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0930_
timestamp 1618216021
transform 1 0 2484 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1618216021
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1618216021
transform 1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1618216021
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1618216021
transform 1 0 2116 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1618216021
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1618216021
transform 1 0 3128 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_28
timestamp 1618216021
transform 1 0 3680 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1618216021
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1618216021
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _0621_
timestamp 1618216021
transform 1 0 6624 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_54
timestamp 1618216021
transform 1 0 6072 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0620_
timestamp 1618216021
transform 1 0 8372 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1618216021
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1618216021
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_78
timestamp 1618216021
transform 1 0 8280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_82
timestamp 1618216021
transform 1 0 8648 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_87
timestamp 1618216021
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1618216021
transform 1 0 10488 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0709_
timestamp 1618216021
transform 1 0 9476 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1618216021
transform 1 0 11132 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_97
timestamp 1618216021
transform 1 0 10028 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1618216021
transform 1 0 10396 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_105
timestamp 1618216021
transform 1 0 10764 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_2  _0711_
timestamp 1618216021
transform 1 0 12972 0 -1 23392
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_38_125
timestamp 1618216021
transform 1 0 12604 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0879_
timestamp 1618216021
transform 1 0 14720 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1618216021
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_139
timestamp 1618216021
transform 1 0 13892 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_144
timestamp 1618216021
transform 1 0 14352 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_152
timestamp 1618216021
transform 1 0 15088 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0729_
timestamp 1618216021
transform 1 0 16008 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_38_160
timestamp 1618216021
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1618216021
transform 1 0 16836 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0976_
timestamp 1618216021
transform 1 0 17848 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_i_clk
timestamp 1618216021
transform 1 0 18860 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_i_clk
timestamp 1618216021
transform 1 0 17204 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_178
timestamp 1618216021
transform 1 0 17480 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_189
timestamp 1618216021
transform 1 0 18492 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_196
timestamp 1618216021
transform 1 0 19136 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0877_
timestamp 1618216021
transform 1 0 20056 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1618216021
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_201
timestamp 1618216021
transform 1 0 19596 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_205
timestamp 1618216021
transform 1 0 19964 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_213
timestamp 1618216021
transform 1 0 20700 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1618216021
transform 1 0 21528 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_221
timestamp 1618216021
transform 1 0 21436 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1618216021
transform 1 0 23000 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1618216021
transform 1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1618216021
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_i_clk
timestamp 1618216021
transform 1 0 24012 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_245
timestamp 1618216021
transform 1 0 23644 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_252
timestamp 1618216021
transform 1 0 24288 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_256
timestamp 1618216021
transform 1 0 24656 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1618216021
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1618216021
transform 1 0 26036 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_270
timestamp 1618216021
transform 1 0 25944 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1618216021
transform -1 0 28428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_287
timestamp 1618216021
transform 1 0 27508 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_293
timestamp 1618216021
transform 1 0 28060 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1024_
timestamp 1618216021
transform 1 0 1748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1618216021
transform 1 0 2484 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1618216021
transform 1 0 1932 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1618216021
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1618216021
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1618216021
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1618216021
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1618216021
transform 1 0 1380 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1618216021
transform 1 0 4784 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0932_
timestamp 1618216021
transform 1 0 4232 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1618216021
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_31
timestamp 1618216021
transform 1 0 3956 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_39
timestamp 1618216021
transform 1 0 4692 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_43
timestamp 1618216021
transform 1 0 5060 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_25
timestamp 1618216021
transform 1 0 3404 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_30
timestamp 1618216021
transform 1 0 3864 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_41
timestamp 1618216021
transform 1 0 4876 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0643_
timestamp 1618216021
transform 1 0 5428 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0926_
timestamp 1618216021
transform 1 0 5244 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1618216021
transform 1 0 6072 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1618216021
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_53
timestamp 1618216021
transform 1 0 5980 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1618216021
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_49
timestamp 1618216021
transform 1 0 5612 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_53
timestamp 1618216021
transform 1 0 5980 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0912_
timestamp 1618216021
transform 1 0 7544 0 1 23392
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0916_
timestamp 1618216021
transform 1 0 8004 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1618216021
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_80
timestamp 1618216021
transform 1 0 8464 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1618216021
transform 1 0 7544 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_74
timestamp 1618216021
transform 1 0 7912 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_82
timestamp 1618216021
transform 1 0 8648 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_87
timestamp 1618216021
transform 1 0 9108 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0710_
timestamp 1618216021
transform 1 0 10396 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0981_
timestamp 1618216021
transform 1 0 9384 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1618216021
transform 1 0 9844 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_39_88
timestamp 1618216021
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1618216021
transform 1 0 10028 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1618216021
transform 1 0 13064 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0882_
timestamp 1618216021
transform 1 0 13064 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1618216021
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_110
timestamp 1618216021
transform 1 0 11224 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1618216021
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_127
timestamp 1618216021
transform 1 0 12788 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1618216021
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_123
timestamp 1618216021
transform 1 0 12420 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_129
timestamp 1618216021
transform 1 0 12972 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1618216021
transform 1 0 14076 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0881_
timestamp 1618216021
transform 1 0 14720 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1618216021
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_137
timestamp 1618216021
transform 1 0 13708 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_144
timestamp 1618216021
transform 1 0 14352 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_152
timestamp 1618216021
transform 1 0 15088 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_133
timestamp 1618216021
transform 1 0 13340 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1618216021
transform 1 0 14076 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_144
timestamp 1618216021
transform 1 0 14352 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1618216021
transform 1 0 15732 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0977_
timestamp 1618216021
transform 1 0 15180 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0978_
timestamp 1618216021
transform 1 0 15916 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1618216021
transform 1 0 15548 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1618216021
transform 1 0 15364 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1618216021
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_165
timestamp 1618216021
transform 1 0 16284 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1618216021
transform 1 0 16928 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_174
timestamp 1618216021
transform 1 0 17112 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_162
timestamp 1618216021
transform 1 0 16008 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0919_
timestamp 1618216021
transform 1 0 17296 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0920_
timestamp 1618216021
transform 1 0 17388 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1618216021
transform 1 0 18124 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1618216021
transform 1 0 17664 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_184
timestamp 1618216021
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_181
timestamp 1618216021
transform 1 0 17756 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_193
timestamp 1618216021
transform 1 0 18860 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1618216021
transform 1 0 20516 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1618216021
transform 1 0 20056 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1618216021
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1618216021
transform 1 0 19688 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_199
timestamp 1618216021
transform 1 0 19412 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_201
timestamp 1618216021
transform 1 0 19596 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_209
timestamp 1618216021
transform 1 0 20332 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_214
timestamp 1618216021
transform 1 0 20792 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_218
timestamp 1618216021
transform 1 0 21160 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0678_
timestamp 1618216021
transform 1 0 22540 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0685_
timestamp 1618216021
transform 1 0 22724 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _0686_
timestamp 1618216021
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1618216021
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_222
timestamp 1618216021
transform 1 0 21528 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_229
timestamp 1618216021
transform 1 0 22172 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_240
timestamp 1618216021
transform 1 0 23184 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_231
timestamp 1618216021
transform 1 0 22356 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1200_
timestamp 1618216021
transform 1 0 23920 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1618216021
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_242
timestamp 1618216021
transform 1 0 23368 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_254
timestamp 1618216021
transform 1 0 24472 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_258
timestamp 1618216021
transform 1 0 24840 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1618216021
transform 1 0 25392 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0923_
timestamp 1618216021
transform 1 0 26128 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1618216021
transform 1 0 26036 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_39_264
timestamp 1618216021
transform 1 0 25392 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_279
timestamp 1618216021
transform 1 0 26772 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_267
timestamp 1618216021
transform 1 0 25668 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1618216021
transform -1 0 28428 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1618216021
transform -1 0 28428 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1618216021
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_286
timestamp 1618216021
transform 1 0 27416 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_287
timestamp 1618216021
transform 1 0 27508 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1618216021
transform 1 0 28060 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0928_
timestamp 1618216021
transform 1 0 2208 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1618216021
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1618216021
transform 1 0 1472 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_3
timestamp 1618216021
transform 1 0 1380 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_8
timestamp 1618216021
transform 1 0 1840 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1618216021
transform 1 0 2852 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0927_
timestamp 1618216021
transform 1 0 5060 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1618216021
transform 1 0 3220 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_39
timestamp 1618216021
transform 1 0 4692 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0913_
timestamp 1618216021
transform 1 0 6900 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1618216021
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1618216021
transform 1 0 5428 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_55
timestamp 1618216021
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_58
timestamp 1618216021
transform 1 0 6440 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_62
timestamp 1618216021
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1618216021
transform 1 0 7636 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_67
timestamp 1618216021
transform 1 0 7268 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_87
timestamp 1618216021
transform 1 0 9108 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0717_
timestamp 1618216021
transform 1 0 10028 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_41_95
timestamp 1618216021
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1618216021
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1618216021
transform 1 0 12052 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _0718_
timestamp 1618216021
transform 1 0 12696 0 1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1618216021
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1618216021
transform 1 0 11684 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_122
timestamp 1618216021
transform 1 0 12328 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0692_
timestamp 1618216021
transform 1 0 13984 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0701_
timestamp 1618216021
transform 1 0 15088 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_41_136
timestamp 1618216021
transform 1 0 13616 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1618216021
transform 1 0 14628 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_151
timestamp 1618216021
transform 1 0 14996 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1618216021
transform 1 0 16192 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1618216021
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_159
timestamp 1618216021
transform 1 0 15732 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_163
timestamp 1618216021
transform 1 0 16100 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_167
timestamp 1618216021
transform 1 0 16468 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1618216021
transform 1 0 16928 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0702_
timestamp 1618216021
transform 1 0 17296 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1618216021
transform 1 0 18768 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1618216021
transform 1 0 18400 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_195
timestamp 1618216021
transform 1 0 19044 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1618216021
transform 1 0 21160 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_207
timestamp 1618216021
transform 1 0 20148 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_215
timestamp 1618216021
transform 1 0 20884 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1618216021
transform 1 0 23000 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1618216021
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_221
timestamp 1618216021
transform 1 0 21436 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_227
timestamp 1618216021
transform 1 0 21988 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_229
timestamp 1618216021
transform 1 0 22172 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_237
timestamp 1618216021
transform 1 0 22908 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1618216021
transform 1 0 24012 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_245
timestamp 1618216021
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0925_
timestamp 1618216021
transform 1 0 26128 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_41_265
timestamp 1618216021
transform 1 0 25484 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_271
timestamp 1618216021
transform 1 0 26036 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_279
timestamp 1618216021
transform 1 0 26772 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1618216021
transform -1 0 28428 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1618216021
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_286
timestamp 1618216021
transform 1 0 27416 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0931_
timestamp 1618216021
transform 1 0 2760 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1618216021
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1618216021
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_6
timestamp 1618216021
transform 1 0 1656 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1618216021
transform 1 0 4232 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1618216021
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_25
timestamp 1618216021
transform 1 0 3404 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_30
timestamp 1618216021
transform 1 0 3864 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_37
timestamp 1618216021
transform 1 0 4508 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_43
timestamp 1618216021
transform 1 0 5060 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0918_
timestamp 1618216021
transform 1 0 7084 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1618216021
transform 1 0 5152 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_60
timestamp 1618216021
transform 1 0 6624 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_64
timestamp 1618216021
transform 1 0 6992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _0716_
timestamp 1618216021
transform 1 0 8096 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1618216021
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_72
timestamp 1618216021
transform 1 0 7728 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_82
timestamp 1618216021
transform 1 0 8648 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_87
timestamp 1618216021
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1618216021
transform 1 0 10120 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1618216021
transform 1 0 9476 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0835_
timestamp 1618216021
transform 1 0 10856 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_42_94
timestamp 1618216021
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1618216021
transform 1 0 10396 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1618216021
transform 1 0 10764 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0880_
timestamp 1618216021
transform 1 0 12236 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_42_113
timestamp 1618216021
transform 1 0 11500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1618216021
transform 1 0 12880 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1618216021
transform 1 0 13248 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1618216021
transform 1 0 14720 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1618216021
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_139
timestamp 1618216021
transform 1 0 13892 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_144
timestamp 1618216021
transform 1 0 14352 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1618216021
transform 1 0 16652 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_164
timestamp 1618216021
transform 1 0 16192 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_168
timestamp 1618216021
transform 1 0 16560 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_172
timestamp 1618216021
transform 1 0 16928 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1618216021
transform 1 0 18768 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_2  _0730_
timestamp 1618216021
transform 1 0 17296 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_188
timestamp 1618216021
transform 1 0 18400 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_195
timestamp 1618216021
transform 1 0 19044 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1618216021
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_199
timestamp 1618216021
transform 1 0 19412 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1618216021
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1618216021
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0687_
timestamp 1618216021
transform 1 0 22816 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1618216021
transform 1 0 21804 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_233
timestamp 1618216021
transform 1 0 22540 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1618216021
transform 1 0 25208 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1618216021
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_243
timestamp 1618216021
transform 1 0 23460 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_255
timestamp 1618216021
transform 1 0 24564 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1618216021
transform 1 0 24840 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1044_
timestamp 1618216021
transform 1 0 27048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_278
timestamp 1618216021
transform 1 0 26680 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1618216021
transform -1 0 28428 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_286
timestamp 1618216021
transform 1 0 27416 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1023_
timestamp 1618216021
transform 1 0 2116 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1618216021
transform 1 0 2852 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1618216021
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1618216021
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1618216021
transform 1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_15
timestamp 1618216021
transform 1 0 2484 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_35
timestamp 1618216021
transform 1 0 4324 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_43
timestamp 1618216021
transform 1 0 5060 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _0636_
timestamp 1618216021
transform 1 0 6808 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0929_
timestamp 1618216021
transform 1 0 5244 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1618216021
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1618216021
transform 1 0 5888 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_56
timestamp 1618216021
transform 1 0 6256 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_58
timestamp 1618216021
transform 1 0 6440 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1618216021
transform 1 0 7728 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_68
timestamp 1618216021
transform 1 0 7360 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_75
timestamp 1618216021
transform 1 0 8004 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_87
timestamp 1618216021
transform 1 0 9108 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1618216021
transform 1 0 9752 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_43_93
timestamp 1618216021
transform 1 0 9660 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0832_
timestamp 1618216021
transform 1 0 12052 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1618216021
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_110
timestamp 1618216021
transform 1 0 11224 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_115
timestamp 1618216021
transform 1 0 11684 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_126
timestamp 1618216021
transform 1 0 12696 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _0693_
timestamp 1618216021
transform 1 0 13248 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _0836_
timestamp 1618216021
transform 1 0 15824 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1618216021
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_153
timestamp 1618216021
transform 1 0 15180 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_159
timestamp 1618216021
transform 1 0 15732 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_167
timestamp 1618216021
transform 1 0 16468 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_172
timestamp 1618216021
transform 1 0 16928 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1618216021
transform 1 0 17296 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_43_192
timestamp 1618216021
transform 1 0 18768 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0719_
timestamp 1618216021
transform 1 0 20884 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_43_204
timestamp 1618216021
transform 1 0 19872 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_212
timestamp 1618216021
transform 1 0 20608 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1618216021
transform 1 0 22816 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1618216021
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_222
timestamp 1618216021
transform 1 0 21528 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_229
timestamp 1618216021
transform 1 0 22172 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_235
timestamp 1618216021
transform 1 0 22724 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0694_
timestamp 1618216021
transform 1 0 24656 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1618216021
transform 1 0 24288 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1618216021
transform 1 0 26588 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_263
timestamp 1618216021
transform 1 0 25300 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_275
timestamp 1618216021
transform 1 0 26404 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1618216021
transform 1 0 26956 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1618216021
transform -1 0 28428 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1618216021
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_286
timestamp 1618216021
transform 1 0 27416 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1618216021
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1618216021
transform 1 0 1748 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1618216021
transform 1 0 1380 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_11
timestamp 1618216021
transform 1 0 2116 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1618216021
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_23
timestamp 1618216021
transform 1 0 3220 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_30
timestamp 1618216021
transform 1 0 3864 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_42
timestamp 1618216021
transform 1 0 4968 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_54
timestamp 1618216021
transform 1 0 6072 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1618216021
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1618216021
transform 1 0 7176 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_78
timestamp 1618216021
transform 1 0 8280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_87
timestamp 1618216021
transform 1 0 9108 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1618216021
transform 1 0 9476 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_44_107
timestamp 1618216021
transform 1 0 10948 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1618216021
transform 1 0 11776 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_44_115
timestamp 1618216021
transform 1 0 11684 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1618216021
transform 1 0 13616 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1618216021
transform 1 0 15088 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1618216021
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_132
timestamp 1618216021
transform 1 0 13248 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_139
timestamp 1618216021
transform 1 0 13892 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1618216021
transform 1 0 14352 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1618216021
transform 1 0 17112 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_44_168
timestamp 1618216021
transform 1 0 16560 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_190
timestamp 1618216021
transform 1 0 18584 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1618216021
transform 1 0 20884 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1618216021
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_198
timestamp 1618216021
transform 1 0 19320 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1618216021
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_213
timestamp 1618216021
transform 1 0 20700 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1618216021
transform 1 0 22908 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_44_231
timestamp 1618216021
transform 1 0 22356 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1618216021
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1618216021
transform 1 0 24380 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1618216021
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1618216021
transform 1 0 26680 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_270
timestamp 1618216021
transform 1 0 25944 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_282
timestamp 1618216021
transform 1 0 27048 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1618216021
transform -1 0 28428 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1618216021
transform 1 0 27416 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_290
timestamp 1618216021
transform 1 0 27784 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1618216021
transform 1 0 2116 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1618216021
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 1618216021
transform 1 0 1380 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1618216021
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1618216021
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1618216021
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0917_
timestamp 1618216021
transform 1 0 7084 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1618216021
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_51
timestamp 1618216021
transform 1 0 5796 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_58
timestamp 1618216021
transform 1 0 6440 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_64
timestamp 1618216021
transform 1 0 6992 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1618216021
transform 1 0 8096 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_72
timestamp 1618216021
transform 1 0 7728 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_83
timestamp 1618216021
transform 1 0 8740 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0982_
timestamp 1618216021
transform 1 0 9568 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1618216021
transform 1 0 10580 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_91
timestamp 1618216021
transform 1 0 9476 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1618216021
transform 1 0 10212 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1618216021
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1618216021
transform 1 0 12052 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1618216021
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1618216021
transform 1 0 11684 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1618216021
transform 1 0 13892 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1618216021
transform 1 0 14996 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_135
timestamp 1618216021
transform 1 0 13524 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_142
timestamp 1618216021
transform 1 0 14168 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_150
timestamp 1618216021
transform 1 0 14904 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1618216021
transform 1 0 16100 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1618216021
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_158
timestamp 1618216021
transform 1 0 15640 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_162
timestamp 1618216021
transform 1 0 16008 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_166
timestamp 1618216021
transform 1 0 16376 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_170
timestamp 1618216021
transform 1 0 16744 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1618216021
transform 1 0 16928 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1618216021
transform 1 0 18308 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1618216021
transform 1 0 18952 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1618216021
transform 1 0 17296 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_183
timestamp 1618216021
transform 1 0 17940 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1618216021
transform 1 0 18584 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_197
timestamp 1618216021
transform 1 0 19228 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_209
timestamp 1618216021
transform 1 0 20332 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1618216021
transform 1 0 21436 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1618216021
transform 1 0 22816 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1618216021
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_224
timestamp 1618216021
transform 1 0 21712 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_229
timestamp 1618216021
transform 1 0 22172 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_235
timestamp 1618216021
transform 1 0 22724 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_243
timestamp 1618216021
transform 1 0 23460 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_255
timestamp 1618216021
transform 1 0 24564 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output159
timestamp 1618216021
transform 1 0 26588 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_267
timestamp 1618216021
transform 1 0 25668 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_275
timestamp 1618216021
transform 1 0 26404 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1618216021
transform 1 0 26956 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1618216021
transform -1 0 28428 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1618216021
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_286
timestamp 1618216021
transform 1 0 27416 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1618216021
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1618216021
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1618216021
transform 1 0 1380 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1618216021
transform 1 0 1748 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1618216021
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_6
timestamp 1618216021
transform 1 0 1656 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_10
timestamp 1618216021
transform 1 0 2024 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1618216021
transform 1 0 2116 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1618216021
transform 1 0 2760 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_14
timestamp 1618216021
transform 1 0 2392 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_21
timestamp 1618216021
transform 1 0 3036 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_10
timestamp 1618216021
transform 1 0 2024 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1618216021
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1618216021
transform 1 0 3404 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1618216021
transform 1 0 3128 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_28
timestamp 1618216021
transform 1 0 3680 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1618216021
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1618216021
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_28
timestamp 1618216021
transform 1 0 3680 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_40
timestamp 1618216021
transform 1 0 4784 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1618216021
transform 1 0 6348 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1618216021
transform 1 0 6808 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1618216021
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_54
timestamp 1618216021
transform 1 0 6072 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1618216021
transform 1 0 5888 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_56
timestamp 1618216021
transform 1 0 6256 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_58
timestamp 1618216021
transform 1 0 6440 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1618216021
transform 1 0 8648 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1618216021
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1618216021
transform 1 0 8188 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1618216021
transform 1 0 7820 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_80
timestamp 1618216021
transform 1 0 8464 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_87
timestamp 1618216021
transform 1 0 9108 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_78
timestamp 1618216021
transform 1 0 8280 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1618216021
transform 1 0 9476 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0979_
timestamp 1618216021
transform 1 0 10120 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1036_
timestamp 1618216021
transform 1 0 10488 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_94
timestamp 1618216021
transform 1 0 9752 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1618216021
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_98
timestamp 1618216021
transform 1 0 10120 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1618216021
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1618216021
transform 1 0 11868 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1618216021
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1618216021
transform 1 0 12052 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_115
timestamp 1618216021
transform 1 0 11684 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_122
timestamp 1618216021
transform 1 0 12328 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0980_
timestamp 1618216021
transform 1 0 14720 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1618216021
transform 1 0 14352 0 1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1618216021
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1618216021
transform 1 0 13708 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_133
timestamp 1618216021
transform 1 0 13340 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1618216021
transform 1 0 14076 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_144
timestamp 1618216021
transform 1 0 14352 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_134
timestamp 1618216021
transform 1 0 13432 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1618216021
transform 1 0 13984 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0983_
timestamp 1618216021
transform 1 0 15732 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1618216021
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1618216021
transform 1 0 16744 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_155
timestamp 1618216021
transform 1 0 15364 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1618216021
transform 1 0 16376 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_173
timestamp 1618216021
transform 1 0 17020 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_161
timestamp 1618216021
transform 1 0 15916 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1618216021
transform 1 0 16652 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_172
timestamp 1618216021
transform 1 0 16928 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0921_
timestamp 1618216021
transform 1 0 17480 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1618216021
transform 1 0 17480 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1618216021
transform 1 0 18492 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_177
timestamp 1618216021
transform 1 0 17388 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1618216021
transform 1 0 18124 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1618216021
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1618216021
transform 1 0 18952 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0924_
timestamp 1618216021
transform 1 0 20240 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1016_
timestamp 1618216021
transform 1 0 19320 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1618216021
transform 1 0 20332 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1618216021
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_201
timestamp 1618216021
transform 1 0 19596 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_202
timestamp 1618216021
transform 1 0 19688 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_215
timestamp 1618216021
transform 1 0 20884 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1020_
timestamp 1618216021
transform 1 0 21252 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1618216021
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1618216021
transform 1 0 22540 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1618216021
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1618216021
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_223
timestamp 1618216021
transform 1 0 21620 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_227
timestamp 1618216021
transform 1 0 21988 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_229
timestamp 1618216021
transform 1 0 22172 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_236
timestamp 1618216021
transform 1 0 22816 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1029_
timestamp 1618216021
transform 1 0 24564 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1618216021
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1618216021
transform 1 0 23920 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_249
timestamp 1618216021
transform 1 0 24012 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_258
timestamp 1618216021
transform 1 0 24840 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1618216021
transform 1 0 24196 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_259
timestamp 1618216021
transform 1 0 24932 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1618216021
transform 1 0 25300 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output158
timestamp 1618216021
transform 1 0 25484 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_264
timestamp 1618216021
transform 1 0 25392 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_266
timestamp 1618216021
transform 1 0 25576 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1018_
timestamp 1618216021
transform 1 0 25944 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_269
timestamp 1618216021
transform 1 0 25852 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output156
timestamp 1618216021
transform 1 0 26220 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_274
timestamp 1618216021
transform 1 0 26312 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1047_
timestamp 1618216021
transform 1 0 26956 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1618216021
transform 1 0 26680 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_277
timestamp 1618216021
transform 1 0 26588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1618216021
transform 1 0 26956 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1618216021
transform -1 0 28428 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1618216021
transform -1 0 28428 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1618216021
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_285
timestamp 1618216021
transform 1 0 27324 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_293
timestamp 1618216021
transform 1 0 28060 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_286
timestamp 1618216021
transform 1 0 27416 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1618216021
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1618216021
transform 1 0 2852 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output154
timestamp 1618216021
transform 1 0 1748 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1618216021
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_11
timestamp 1618216021
transform 1 0 2116 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1618216021
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1618216021
transform 1 0 5060 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1618216021
transform 1 0 4232 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_23
timestamp 1618216021
transform 1 0 3220 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_30
timestamp 1618216021
transform 1 0 3864 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_37
timestamp 1618216021
transform 1 0 4508 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1030_
timestamp 1618216021
transform 1 0 6164 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_46
timestamp 1618216021
transform 1 0 5336 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_54
timestamp 1618216021
transform 1 0 6072 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_59
timestamp 1618216021
transform 1 0 6532 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0915_
timestamp 1618216021
transform 1 0 7268 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1618216021
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1618216021
transform 1 0 8280 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_74
timestamp 1618216021
transform 1 0 7912 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_81
timestamp 1618216021
transform 1 0 8556 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_85
timestamp 1618216021
transform 1 0 8924 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_87
timestamp 1618216021
transform 1 0 9108 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1022_
timestamp 1618216021
transform 1 0 9476 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1618216021
transform 1 0 10212 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_95
timestamp 1618216021
transform 1 0 9844 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1618216021
transform 1 0 12052 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1618216021
transform 1 0 12696 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_115
timestamp 1618216021
transform 1 0 11684 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_122
timestamp 1618216021
transform 1 0 12328 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_129
timestamp 1618216021
transform 1 0 12972 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1618216021
transform 1 0 14720 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1618216021
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1618216021
transform 1 0 13340 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_136
timestamp 1618216021
transform 1 0 13616 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_142
timestamp 1618216021
transform 1 0 14168 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_144
timestamp 1618216021
transform 1 0 14352 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1618216021
transform 1 0 16560 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_164
timestamp 1618216021
transform 1 0 16192 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_171
timestamp 1618216021
transform 1 0 16836 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1618216021
transform 1 0 17480 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_177
timestamp 1618216021
transform 1 0 17388 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_194
timestamp 1618216021
transform 1 0 18952 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1021_
timestamp 1618216021
transform 1 0 20056 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1034_
timestamp 1618216021
transform 1 0 20792 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1618216021
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_201
timestamp 1618216021
transform 1 0 19596 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_205
timestamp 1618216021
transform 1 0 19964 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1618216021
transform 1 0 20424 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_218
timestamp 1618216021
transform 1 0 21160 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1041_
timestamp 1618216021
transform 1 0 21528 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1618216021
transform 1 0 22264 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_226
timestamp 1618216021
transform 1 0 21896 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_233
timestamp 1618216021
transform 1 0 22540 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1618216021
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1618216021
transform 1 0 23368 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1618216021
transform 1 0 24012 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_241
timestamp 1618216021
transform 1 0 23276 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_245
timestamp 1618216021
transform 1 0 23644 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1618216021
transform 1 0 24380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_258
timestamp 1618216021
transform 1 0 24840 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1019_
timestamp 1618216021
transform 1 0 26956 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1618216021
transform 1 0 26220 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1618216021
transform 1 0 25484 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_264
timestamp 1618216021
transform 1 0 25392 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_269
timestamp 1618216021
transform 1 0 25852 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_277
timestamp 1618216021
transform 1 0 26588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1618216021
transform -1 0 28428 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_285
timestamp 1618216021
transform 1 0 27324 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_293
timestamp 1618216021
transform 1 0 28060 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1618216021
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1618216021
transform 1 0 1748 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1618216021
transform 1 0 2484 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1618216021
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1618216021
transform 1 0 2116 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_19
timestamp 1618216021
transform 1 0 2852 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1618216021
transform 1 0 3772 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output149
timestamp 1618216021
transform 1 0 4232 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_27
timestamp 1618216021
transform 1 0 3588 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_30
timestamp 1618216021
transform 1 0 3864 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_38
timestamp 1618216021
transform 1 0 4600 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1618216021
transform 1 0 6440 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1618216021
transform 1 0 5520 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1618216021
transform 1 0 6900 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_46
timestamp 1618216021
transform 1 0 5336 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_52
timestamp 1618216021
transform 1 0 5888 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_59
timestamp 1618216021
transform 1 0 6532 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1618216021
transform 1 0 9108 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1618216021
transform 1 0 8372 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1618216021
transform 1 0 7636 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_67
timestamp 1618216021
transform 1 0 7268 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_75
timestamp 1618216021
transform 1 0 8004 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_83
timestamp 1618216021
transform 1 0 8740 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1618216021
transform 1 0 10580 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1618216021
transform 1 0 9844 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_88
timestamp 1618216021
transform 1 0 9200 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_94
timestamp 1618216021
transform 1 0 9752 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1618216021
transform 1 0 10212 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_107
timestamp 1618216021
transform 1 0 10948 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1618216021
transform 1 0 11776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1618216021
transform 1 0 12420 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1618216021
transform 1 0 13156 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_115
timestamp 1618216021
transform 1 0 11684 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_117
timestamp 1618216021
transform 1 0 11868 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_127
timestamp 1618216021
transform 1 0 12788 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1618216021
transform 1 0 14444 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1618216021
transform 1 0 14904 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1618216021
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_143
timestamp 1618216021
transform 1 0 14260 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1618216021
transform 1 0 14536 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1618216021
transform 1 0 17112 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1618216021
transform 1 0 16376 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1618216021
transform 1 0 15640 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1618216021
transform 1 0 15272 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_162
timestamp 1618216021
transform 1 0 16008 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_170
timestamp 1618216021
transform 1 0 16744 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1618216021
transform 1 0 17572 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1618216021
transform 1 0 18584 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_175
timestamp 1618216021
transform 1 0 17204 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_186
timestamp 1618216021
transform 1 0 18216 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_194
timestamp 1618216021
transform 1 0 18952 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1618216021
transform 1 0 19780 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1618216021
transform 1 0 20700 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_202
timestamp 1618216021
transform 1 0 19688 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_204
timestamp 1618216021
transform 1 0 19872 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_212
timestamp 1618216021
transform 1 0 20608 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1618216021
transform 1 0 21068 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1618216021
transform 1 0 22448 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1618216021
transform 1 0 21620 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1618216021
transform 1 0 22908 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_227
timestamp 1618216021
transform 1 0 21988 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1618216021
transform 1 0 22356 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_233
timestamp 1618216021
transform 1 0 22540 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1618216021
transform 1 0 25116 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1618216021
transform 1 0 23644 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1618216021
transform 1 0 24380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_241
timestamp 1618216021
transform 1 0 23276 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_249
timestamp 1618216021
transform 1 0 24012 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_257
timestamp 1618216021
transform 1 0 24748 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1618216021
transform 1 0 25208 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1618216021
transform 1 0 27048 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1618216021
transform 1 0 26312 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1618216021
transform 1 0 25576 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_270
timestamp 1618216021
transform 1 0 25944 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_278
timestamp 1618216021
transform 1 0 26680 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1618216021
transform -1 0 28428 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1618216021
transform 1 0 27784 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1618216021
transform 1 0 27416 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_291
timestamp 1618216021
transform 1 0 27876 0 1 28832
box -38 -48 314 592
<< labels >>
rlabel metal3 s 28780 22448 29580 22568 4 i_clk
port 1 nsew
rlabel metal3 s 0 27888 800 28008 4 i_copro_crm[0]
port 2 nsew
rlabel metal3 s 0 12928 800 13048 4 i_copro_crm[1]
port 3 nsew
rlabel metal2 s 13358 0 13414 800 4 i_copro_crm[2]
port 4 nsew
rlabel metal2 s 25318 30924 25374 31724 4 i_copro_crm[3]
port 5 nsew
rlabel metal2 s 6918 30924 6974 31724 4 i_copro_crn[0]
port 6 nsew
rlabel metal2 s 17038 30924 17094 31724 4 i_copro_crn[1]
port 7 nsew
rlabel metal2 s 5998 0 6054 800 4 i_copro_crn[2]
port 8 nsew
rlabel metal3 s 0 29248 800 29368 4 i_copro_crn[3]
port 9 nsew
rlabel metal2 s 16118 30924 16174 31724 4 i_copro_num[0]
port 10 nsew
rlabel metal3 s 28780 9528 29580 9648 4 i_copro_num[1]
port 11 nsew
rlabel metal2 s 26238 30924 26294 31724 4 i_copro_num[2]
port 12 nsew
rlabel metal2 s 17038 0 17094 800 4 i_copro_num[3]
port 13 nsew
rlabel metal2 s 9678 30924 9734 31724 4 i_copro_opcode1[0]
port 14 nsew
rlabel metal3 s 0 8848 800 8968 4 i_copro_opcode1[1]
port 15 nsew
rlabel metal2 s 21178 0 21234 800 4 i_copro_opcode1[2]
port 16 nsew
rlabel metal2 s 7378 30924 7434 31724 4 i_copro_opcode2[0]
port 17 nsew
rlabel metal2 s 13358 30924 13414 31724 4 i_copro_opcode2[1]
port 18 nsew
rlabel metal2 s 6918 0 6974 800 4 i_copro_opcode2[2]
port 19 nsew
rlabel metal3 s 0 23128 800 23248 4 i_copro_operation[0]
port 20 nsew
rlabel metal3 s 0 25168 800 25288 4 i_copro_operation[1]
port 21 nsew
rlabel metal2 s 1858 30924 1914 31724 4 i_copro_write_data[0]
port 22 nsew
rlabel metal2 s 20258 30924 20314 31724 4 i_copro_write_data[10]
port 23 nsew
rlabel metal2 s 5078 30924 5134 31724 4 i_copro_write_data[11]
port 24 nsew
rlabel metal2 s 17498 0 17554 800 4 i_copro_write_data[12]
port 25 nsew
rlabel metal3 s 28780 6808 29580 6928 4 i_copro_write_data[13]
port 26 nsew
rlabel metal2 s 23478 30924 23534 31724 4 i_copro_write_data[14]
port 27 nsew
rlabel metal2 s 5078 0 5134 800 4 i_copro_write_data[15]
port 28 nsew
rlabel metal2 s 28538 0 28594 800 4 i_copro_write_data[16]
port 29 nsew
rlabel metal2 s 4618 0 4674 800 4 i_copro_write_data[17]
port 30 nsew
rlabel metal2 s 18878 0 18934 800 4 i_copro_write_data[18]
port 31 nsew
rlabel metal3 s 28780 23808 29580 23928 4 i_copro_write_data[19]
port 32 nsew
rlabel metal2 s 14738 30924 14794 31724 4 i_copro_write_data[1]
port 33 nsew
rlabel metal2 s 12438 30924 12494 31724 4 i_copro_write_data[20]
port 34 nsew
rlabel metal2 s 21638 30924 21694 31724 4 i_copro_write_data[21]
port 35 nsew
rlabel metal3 s 0 9528 800 9648 4 i_copro_write_data[22]
port 36 nsew
rlabel metal3 s 28780 20408 29580 20528 4 i_copro_write_data[23]
port 37 nsew
rlabel metal3 s 0 6128 800 6248 4 i_copro_write_data[24]
port 38 nsew
rlabel metal2 s 8758 0 8814 800 4 i_copro_write_data[25]
port 39 nsew
rlabel metal3 s 28780 14968 29580 15088 4 i_copro_write_data[26]
port 40 nsew
rlabel metal3 s 28780 19728 29580 19848 4 i_copro_write_data[27]
port 41 nsew
rlabel metal2 s 12898 30924 12954 31724 4 i_copro_write_data[28]
port 42 nsew
rlabel metal3 s 28780 4768 29580 4888 4 i_copro_write_data[29]
port 43 nsew
rlabel metal2 s 14278 0 14334 800 4 i_copro_write_data[2]
port 44 nsew
rlabel metal3 s 0 14968 800 15088 4 i_copro_write_data[30]
port 45 nsew
rlabel metal2 s 6458 0 6514 800 4 i_copro_write_data[31]
port 46 nsew
rlabel metal2 s 13818 0 13874 800 4 i_copro_write_data[3]
port 47 nsew
rlabel metal2 s 11518 0 11574 800 4 i_copro_write_data[4]
port 48 nsew
rlabel metal3 s 28780 4088 29580 4208 4 i_copro_write_data[5]
port 49 nsew
rlabel metal2 s 2778 0 2834 800 4 i_copro_write_data[6]
port 50 nsew
rlabel metal2 s 27158 30924 27214 31724 4 i_copro_write_data[7]
port 51 nsew
rlabel metal3 s 0 1368 800 1488 4 i_copro_write_data[8]
port 52 nsew
rlabel metal3 s 28780 21088 29580 21208 4 i_copro_write_data[9]
port 53 nsew
rlabel metal2 s 478 0 534 800 4 i_core_stall
port 54 nsew
rlabel metal3 s 0 12248 800 12368 4 i_fault
port 55 nsew
rlabel metal3 s 0 17008 800 17128 4 i_fault_address[0]
port 56 nsew
rlabel metal2 s 11518 30924 11574 31724 4 i_fault_address[10]
port 57 nsew
rlabel metal3 s 0 6808 800 6928 4 i_fault_address[11]
port 58 nsew
rlabel metal3 s 28780 1368 29580 1488 4 i_fault_address[12]
port 59 nsew
rlabel metal3 s 0 28568 800 28688 4 i_fault_address[13]
port 60 nsew
rlabel metal3 s 28780 10208 29580 10328 4 i_fault_address[14]
port 61 nsew
rlabel metal2 s 938 30924 994 31724 4 i_fault_address[15]
port 62 nsew
rlabel metal2 s 11058 30924 11114 31724 4 i_fault_address[16]
port 63 nsew
rlabel metal2 s 23018 0 23074 800 4 i_fault_address[17]
port 64 nsew
rlabel metal2 s 15198 30924 15254 31724 4 i_fault_address[18]
port 65 nsew
rlabel metal2 s 20718 0 20774 800 4 i_fault_address[19]
port 66 nsew
rlabel metal2 s 22558 0 22614 800 4 i_fault_address[1]
port 67 nsew
rlabel metal2 s 9218 30924 9274 31724 4 i_fault_address[20]
port 68 nsew
rlabel metal2 s 18418 30924 18474 31724 4 i_fault_address[21]
port 69 nsew
rlabel metal3 s 0 4088 800 4208 4 i_fault_address[22]
port 70 nsew
rlabel metal2 s 4158 0 4214 800 4 i_fault_address[23]
port 71 nsew
rlabel metal3 s 28780 7488 29580 7608 4 i_fault_address[24]
port 72 nsew
rlabel metal3 s 0 15648 800 15768 4 i_fault_address[25]
port 73 nsew
rlabel metal3 s 28780 3408 29580 3528 4 i_fault_address[26]
port 74 nsew
rlabel metal2 s 4158 30924 4214 31724 4 i_fault_address[27]
port 75 nsew
rlabel metal2 s 24858 0 24914 800 4 i_fault_address[28]
port 76 nsew
rlabel metal2 s 19338 0 19394 800 4 i_fault_address[29]
port 77 nsew
rlabel metal2 s 19798 0 19854 800 4 i_fault_address[2]
port 78 nsew
rlabel metal3 s 0 20408 800 20528 4 i_fault_address[30]
port 79 nsew
rlabel metal3 s 28780 30608 29580 30728 4 i_fault_address[31]
port 80 nsew
rlabel metal2 s 16578 30924 16634 31724 4 i_fault_address[3]
port 81 nsew
rlabel metal2 s 2318 0 2374 800 4 i_fault_address[4]
port 82 nsew
rlabel metal2 s 3238 0 3294 800 4 i_fault_address[5]
port 83 nsew
rlabel metal3 s 28780 15648 29580 15768 4 i_fault_address[6]
port 84 nsew
rlabel metal2 s 2778 30924 2834 31724 4 i_fault_address[7]
port 85 nsew
rlabel metal3 s 0 30608 800 30728 4 i_fault_address[8]
port 86 nsew
rlabel metal3 s 0 3408 800 3528 4 i_fault_address[9]
port 87 nsew
rlabel metal2 s 7838 0 7894 800 4 i_fault_status[0]
port 88 nsew
rlabel metal2 s 15198 0 15254 800 4 i_fault_status[1]
port 89 nsew
rlabel metal2 s 22558 30924 22614 31724 4 i_fault_status[2]
port 90 nsew
rlabel metal2 s 23938 30924 23994 31724 4 i_fault_status[3]
port 91 nsew
rlabel metal2 s 24398 0 24454 800 4 i_fault_status[4]
port 92 nsew
rlabel metal2 s 17958 0 18014 800 4 i_fault_status[5]
port 93 nsew
rlabel metal3 s 28780 688 29580 808 4 i_fault_status[6]
port 94 nsew
rlabel metal3 s 0 4768 800 4888 4 i_fault_status[7]
port 95 nsew
rlabel metal3 s 28780 27888 29580 28008 4 o_cache_enable
port 96 nsew
rlabel metal2 s 27618 30924 27674 31724 4 o_cache_flush
port 97 nsew
rlabel metal2 s 28078 0 28134 800 4 o_cacheable_area[0]
port 98 nsew
rlabel metal3 s 0 10208 800 10328 4 o_cacheable_area[10]
port 99 nsew
rlabel metal3 s 0 26528 800 26648 4 o_cacheable_area[11]
port 100 nsew
rlabel metal2 s 938 0 994 800 4 o_cacheable_area[12]
port 101 nsew
rlabel metal3 s 28780 18368 29580 18488 4 o_cacheable_area[13]
port 102 nsew
rlabel metal2 s 17958 30924 18014 31724 4 o_cacheable_area[14]
port 103 nsew
rlabel metal2 s 5538 30924 5594 31724 4 o_cacheable_area[15]
port 104 nsew
rlabel metal3 s 28780 12248 29580 12368 4 o_cacheable_area[16]
port 105 nsew
rlabel metal3 s 0 7488 800 7608 4 o_cacheable_area[17]
port 106 nsew
rlabel metal2 s 1398 0 1454 800 4 o_cacheable_area[18]
port 107 nsew
rlabel metal2 s 20718 30924 20774 31724 4 o_cacheable_area[19]
port 108 nsew
rlabel metal2 s 19798 30924 19854 31724 4 o_cacheable_area[1]
port 109 nsew
rlabel metal3 s 0 2048 800 2168 4 o_cacheable_area[20]
port 110 nsew
rlabel metal2 s 10598 30924 10654 31724 4 o_cacheable_area[21]
port 111 nsew
rlabel metal2 s 10598 0 10654 800 4 o_cacheable_area[22]
port 112 nsew
rlabel metal2 s 16118 0 16174 800 4 o_cacheable_area[23]
port 113 nsew
rlabel metal3 s 0 17688 800 17808 4 o_cacheable_area[24]
port 114 nsew
rlabel metal3 s 0 18368 800 18488 4 o_cacheable_area[25]
port 115 nsew
rlabel metal2 s 22098 30924 22154 31724 4 o_cacheable_area[26]
port 116 nsew
rlabel metal2 s 9678 0 9734 800 4 o_cacheable_area[27]
port 117 nsew
rlabel metal3 s 28780 17688 29580 17808 4 o_cacheable_area[28]
port 118 nsew
rlabel metal3 s 28780 26528 29580 26648 4 o_cacheable_area[29]
port 119 nsew
rlabel metal2 s 8298 0 8354 800 4 o_cacheable_area[2]
port 120 nsew
rlabel metal3 s 28780 14288 29580 14408 4 o_cacheable_area[30]
port 121 nsew
rlabel metal3 s 0 19728 800 19848 4 o_cacheable_area[31]
port 122 nsew
rlabel metal2 s 28078 30924 28134 31724 4 o_cacheable_area[3]
port 123 nsew
rlabel metal2 s 28998 30924 29054 31724 4 o_cacheable_area[4]
port 124 nsew
rlabel metal2 s 18878 30924 18934 31724 4 o_cacheable_area[5]
port 125 nsew
rlabel metal2 s 14278 30924 14334 31724 4 o_cacheable_area[6]
port 126 nsew
rlabel metal2 s 8758 30924 8814 31724 4 o_cacheable_area[7]
port 127 nsew
rlabel metal3 s 0 25848 800 25968 4 o_cacheable_area[8]
port 128 nsew
rlabel metal3 s 0 23808 800 23928 4 o_cacheable_area[9]
port 129 nsew
rlabel metal2 s 11978 0 12034 800 4 o_copro_read_data[0]
port 130 nsew
rlabel metal3 s 28780 11568 29580 11688 4 o_copro_read_data[10]
port 131 nsew
rlabel metal3 s 28780 25848 29580 25968 4 o_copro_read_data[11]
port 132 nsew
rlabel metal2 s 24398 30924 24454 31724 4 o_copro_read_data[12]
port 133 nsew
rlabel metal3 s 0 22448 800 22568 4 o_copro_read_data[13]
port 134 nsew
rlabel metal3 s 28780 17008 29580 17128 4 o_copro_read_data[14]
port 135 nsew
rlabel metal3 s 28780 12928 29580 13048 4 o_copro_read_data[15]
port 136 nsew
rlabel metal2 s 12438 0 12494 800 4 o_copro_read_data[16]
port 137 nsew
rlabel metal2 s 5998 30924 6054 31724 4 o_copro_read_data[17]
port 138 nsew
rlabel metal2 s 23478 0 23534 800 4 o_copro_read_data[18]
port 139 nsew
rlabel metal2 s 26698 0 26754 800 4 o_copro_read_data[19]
port 140 nsew
rlabel metal2 s 26238 0 26294 800 4 o_copro_read_data[1]
port 141 nsew
rlabel metal3 s 28780 6128 29580 6248 4 o_copro_read_data[20]
port 142 nsew
rlabel metal3 s 28780 2048 29580 2168 4 o_copro_read_data[21]
port 143 nsew
rlabel metal2 s 25778 0 25834 800 4 o_copro_read_data[22]
port 144 nsew
rlabel metal3 s 28780 25168 29580 25288 4 o_copro_read_data[23]
port 145 nsew
rlabel metal2 s 2318 30924 2374 31724 4 o_copro_read_data[24]
port 146 nsew
rlabel metal2 s 21638 0 21694 800 4 o_copro_read_data[25]
port 147 nsew
rlabel metal3 s 28780 8848 29580 8968 4 o_copro_read_data[26]
port 148 nsew
rlabel metal2 s 7838 30924 7894 31724 4 o_copro_read_data[27]
port 149 nsew
rlabel metal2 s 3698 30924 3754 31724 4 o_copro_read_data[28]
port 150 nsew
rlabel metal2 s 15658 0 15714 800 4 o_copro_read_data[29]
port 151 nsew
rlabel metal3 s 0 21088 800 21208 4 o_copro_read_data[2]
port 152 nsew
rlabel metal3 s 0 11568 800 11688 4 o_copro_read_data[30]
port 153 nsew
rlabel metal2 s 27618 0 27674 800 4 o_copro_read_data[31]
port 154 nsew
rlabel metal2 s 478 30924 534 31724 4 o_copro_read_data[3]
port 155 nsew
rlabel metal3 s 28780 23128 29580 23248 4 o_copro_read_data[4]
port 156 nsew
rlabel metal3 s 28780 29248 29580 29368 4 o_copro_read_data[5]
port 157 nsew
rlabel metal3 s 0 14288 800 14408 4 o_copro_read_data[6]
port 158 nsew
rlabel metal2 s 25778 30924 25834 31724 4 o_copro_read_data[7]
port 159 nsew
rlabel metal3 s 28780 28568 29580 28688 4 o_copro_read_data[8]
port 160 nsew
rlabel metal2 s 10138 0 10194 800 4 o_copro_read_data[9]
port 161 nsew
rlabel metal4 s 23714 2128 24034 29424 4 VPWR
port 162 nsew
rlabel metal4 s 14606 2128 14926 29424 4 VPWR
port 162 nsew
rlabel metal4 s 5498 2128 5818 29424 4 VPWR
port 162 nsew
rlabel metal5 s 1104 24635 28428 24955 4 VPWR
port 162 nsew
rlabel metal5 s 1104 15568 28428 15888 4 VPWR
port 162 nsew
rlabel metal5 s 1104 6501 28428 6821 4 VPWR
port 162 nsew
rlabel metal4 s 19160 2128 19480 29424 4 VGND
port 163 nsew
rlabel metal4 s 10052 2128 10372 29424 4 VGND
port 163 nsew
rlabel metal5 s 1104 20101 28428 20421 4 VGND
port 163 nsew
rlabel metal5 s 1104 11035 28428 11355 4 VGND
port 163 nsew
<< properties >>
string FIXED_BBOX 0 0 29580 31724
<< end >>
